--------------------------------------------------------------------------------
--               FPAdderDualPath_8_47_8_47_8_47400_DualSubClose
--                            (IntDualSub_50_400)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdderDualPath_8_47_8_47_8_47400_DualSubClose is
   port ( 
-- OL clk : in std_logic;
-- OL     rst : in std_logic;
          X : in  std_logic_vector(49 downto 0);
          Y : in  std_logic_vector(49 downto 0);
          RxMy : out  std_logic_vector(49 downto 0);
          RyMx : out  std_logic_vector(49 downto 0)   );
end entity;

architecture arch of FPAdderDualPath_8_47_8_47_8_47400_DualSubClose is
signal sX0 :  std_logic_vector(49 downto 0);
signal sY0 :  std_logic_vector(49 downto 0);
signal xMy0 :  std_logic_vector(50 downto 0);
signal yMx0 :  std_logic_vector(50 downto 0);
begin
--   process(clk)
--      begin
--         if clk'event and clk = '1' then
--         end if;
--      end process;
   sX0 <= X(49 downto 0);
   sY0 <= Y(49 downto 0);
   xMy0  <= ("0" & sX0) + ("0" & not(sY0)) + '1';
   yMx0 <= ("0" & sY0) + ("0" & not(sX0))+ '1';
   RxMy <= xMy0(49 downto 0);
   RyMx <= yMx0(49 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                FPAdderDualPath_8_47_8_47_8_47400_LZCShifter
--                   (LZCShifter_49_to_49_counting_64_uid4)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdderDualPath_8_47_8_47_8_47400_LZCShifter is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL     rst : in std_logic;
          I : in  std_logic_vector(48 downto 0);
          Count : out  std_logic_vector(5 downto 0);
          O : out  std_logic_vector(48 downto 0)   );
end entity;

architecture arch of FPAdderDualPath_8_47_8_47_8_47400_LZCShifter is
signal level6 :  std_logic_vector(48 downto 0);
signal count5, count5_d1, count5_d2, count5_d3, count5_d4, count5_d5 : std_logic;
signal level5, level5_d1 :  std_logic_vector(48 downto 0);
signal count4, count4_d1, count4_d2, count4_d3, count4_d4 : std_logic;
signal level4, level4_d1 :  std_logic_vector(48 downto 0);
signal count3, count3_d1, count3_d2, count3_d3 : std_logic;
signal level3, level3_d1 :  std_logic_vector(48 downto 0);
signal count2, count2_d1, count2_d2 : std_logic;
signal level2, level2_d1 :  std_logic_vector(48 downto 0);
signal count1, count1_d1 : std_logic;
signal level1, level1_d1 :  std_logic_vector(48 downto 0);
signal count0 : std_logic;
signal level0 :  std_logic_vector(48 downto 0);
signal sCount :  std_logic_vector(5 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
           if(Enable='1') then
            count5_d1 <=  count5;
            count5_d2 <=  count5_d1;
            count5_d3 <=  count5_d2;
            count5_d4 <=  count5_d3;
            count5_d5 <=  count5_d4;
            level5_d1 <=  level5;
            count4_d1 <=  count4;
            count4_d2 <=  count4_d1;
            count4_d3 <=  count4_d2;
            count4_d4 <=  count4_d3;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
            count3_d2 <=  count3_d1;
            count3_d3 <=  count3_d2;
            level3_d1 <=  level3;
            count2_d1 <=  count2;
            count2_d2 <=  count2_d1;
            level2_d1 <=  level2;
            count1_d1 <=  count1;
            level1_d1 <=  level1;
           end if;
         end if;
      end process;
   level6 <= I ;
   count5<= '1' when level6(48 downto 17) = (48 downto 17=>'0') else '0';
   level5<= level6(48 downto 0) when count5='0' else level6(16 downto 0) & (31 downto 0 => '0');

   ----------------Synchro barrier, entering cycle 1----------------
   count4<= '1' when level5_d1(48 downto 33) = (48 downto 33=>'0') else '0';
   level4<= level5_d1(48 downto 0) when count4='0' else level5_d1(32 downto 0) & (15 downto 0 => '0');

   ----------------Synchro barrier, entering cycle 2----------------
   count3<= '1' when level4_d1(48 downto 41) = (48 downto 41=>'0') else '0';
   level3<= level4_d1(48 downto 0) when count3='0' else level4_d1(40 downto 0) & (7 downto 0 => '0');

   ----------------Synchro barrier, entering cycle 3----------------
   count2<= '1' when level3_d1(48 downto 45) = (48 downto 45=>'0') else '0';
   level2<= level3_d1(48 downto 0) when count2='0' else level3_d1(44 downto 0) & (3 downto 0 => '0');

   ----------------Synchro barrier, entering cycle 4----------------
   count1<= '1' when level2_d1(48 downto 47) = (48 downto 47=>'0') else '0';
   level1<= level2_d1(48 downto 0) when count1='0' else level2_d1(46 downto 0) & (1 downto 0 => '0');

   ----------------Synchro barrier, entering cycle 5----------------
   count0<= '1' when level1_d1(48 downto 48) = (48 downto 48=>'0') else '0';
   level0<= level1_d1(48 downto 0) when count0='0' else level1_d1(47 downto 0) & (0 downto 0 => '0');

   O <= level0;
   sCount <= count5_d5 & count4_d4 & count3_d3 & count2_d2 & count1_d1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--               FPAdderDualPath_8_47_8_47_8_47400_RightShifter
--                      (RightShifter_48_by_max_50_uid6)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdderDualPath_8_47_8_47_8_47400_RightShifter is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL     rst : in std_logic;
          X : in  std_logic_vector(47 downto 0);
          S : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(97 downto 0)   );
end entity;

architecture arch of FPAdderDualPath_8_47_8_47_8_47400_RightShifter is
signal level0 :  std_logic_vector(47 downto 0);
signal ps, ps_d1 :  std_logic_vector(5 downto 0);
signal level1 :  std_logic_vector(48 downto 0);
signal level2 :  std_logic_vector(50 downto 0);
signal level3 :  std_logic_vector(54 downto 0);
signal level4, level4_d1 :  std_logic_vector(62 downto 0);
signal level5 :  std_logic_vector(78 downto 0);
signal level6 :  std_logic_vector(110 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
           if(Enable='1') then
            ps_d1 <=  ps;
            level4_d1 <=  level4;
           end if;
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   ----------------Synchro barrier, entering cycle 1----------------
   level5<=  (15 downto 0 => '0') & level4_d1 when ps_d1(4) = '1' else    level4_d1 & (15 downto 0 => '0');
   level6<=  (31 downto 0 => '0') & level5 when ps_d1(5) = '1' else    level5 & (31 downto 0 => '0');
   R <= level6(110 downto 13);
end architecture;

--------------------------------------------------------------------------------
--                FPAdderDualPath_8_47_8_47_8_47400_fracAddFar
--                          (IntAdder_51_f400_uid8)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdderDualPath_8_47_8_47_8_47400_fracAddFar is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL     rst : in std_logic;
          X : in  std_logic_vector(50 downto 0);
          Y : in  std_logic_vector(50 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(50 downto 0);
          Nc : out  std_logic   );
end entity;

architecture arch of FPAdderDualPath_8_47_8_47_8_47400_fracAddFar is
signal s_sum_l0_idx0 :  std_logic_vector(42 downto 0);
signal s_sum_l0_idx1, s_sum_l0_idx1_d1 :  std_logic_vector(9 downto 0);
signal sum_l0_idx0, sum_l0_idx0_d1 :  std_logic_vector(41 downto 0);
signal c_l0_idx0, c_l0_idx0_d1 :  std_logic_vector(0 downto 0);
-- OL signal sum_l0_idx1 :  std_logic_vector(8 downto 0);
-- OL signal c_l0_idx1 :  std_logic_vector(0 downto 0);
signal s_sum_l1_idx1 :  std_logic_vector(9 downto 0);
signal sum_l1_idx1 :  std_logic_vector(8 downto 0);
-- OL signal c_l1_idx1 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
          if(Enable='1') then
            s_sum_l0_idx1_d1 <=  s_sum_l0_idx1;
            sum_l0_idx0_d1 <=  sum_l0_idx0;
            c_l0_idx0_d1 <=  c_l0_idx0;
          end if;
         end if;
      end process;
   --Alternative
   s_sum_l0_idx0 <= ( "0" & X(41 downto 0)) + ( "0" & Y(41 downto 0)) + Cin;
   s_sum_l0_idx1 <= ( "0" & X(50 downto 42)) + ( "0" & Y(50 downto 42));
   sum_l0_idx0 <= s_sum_l0_idx0(41 downto 0);
   c_l0_idx0 <= s_sum_l0_idx0(42 downto 42);
-- OL    sum_l0_idx1 <= s_sum_l0_idx1(8 downto 0);
-- OL    c_l0_idx1 <= s_sum_l0_idx1(9 downto 9);
   ----------------Synchro barrier, entering cycle 1----------------
   s_sum_l1_idx1 <=  s_sum_l0_idx1_d1 + c_l0_idx0_d1(0 downto 0);
   sum_l1_idx1 <= s_sum_l1_idx1(8 downto 0);
-- OL   c_l1_idx1 <= s_sum_l1_idx1(9 downto 9);
   R <= sum_l1_idx1(8 downto 0) & sum_l0_idx0_d1(41 downto 0);

   Nc <= s_sum_l0_idx1_d1(9); 
end architecture;

--------------------------------------------------------------------------------
--              FPAdderDualPath_8_47_8_47_8_47400_finalRoundAdd
--                          (IntAdder_57_f400_uid14)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdderDualPath_8_47_8_47_8_47400_finalRoundAdd is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL     rst : in std_logic;
          X : in  std_logic_vector(56 downto 0);
          Y : in  std_logic_vector(56 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(56 downto 0);
          Nc : out  std_logic   );
end entity;

architecture arch of FPAdderDualPath_8_47_8_47_8_47400_finalRoundAdd is
signal s_sum_l0_idx0 :  std_logic_vector(38 downto 0);
signal s_sum_l0_idx1, s_sum_l0_idx1_d1 :  std_logic_vector(19 downto 0);
signal sum_l0_idx0, sum_l0_idx0_d1 :  std_logic_vector(37 downto 0);
signal c_l0_idx0, c_l0_idx0_d1 :  std_logic_vector(0 downto 0);
-- OL signal sum_l0_idx1 :  std_logic_vector(18 downto 0);
-- OL signal c_l0_idx1 :  std_logic_vector(0 downto 0);
signal s_sum_l1_idx1 :  std_logic_vector(19 downto 0);
signal sum_l1_idx1 :  std_logic_vector(18 downto 0);
-- OL signal c_l1_idx1 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
           if(Enable='1') then
            s_sum_l0_idx1_d1 <=  s_sum_l0_idx1;
            sum_l0_idx0_d1 <=  sum_l0_idx0;
            c_l0_idx0_d1 <=  c_l0_idx0;
            end if;
         end if;
      end process;
   --Alternative
   s_sum_l0_idx0 <= ( "0" & X(37 downto 0)) + ( "0" & Y(37 downto 0)) + Cin;
   s_sum_l0_idx1 <= ( "0" & X(56 downto 38)) + ( "0" & Y(56 downto 38));
   sum_l0_idx0 <= s_sum_l0_idx0(37 downto 0);
   c_l0_idx0 <= s_sum_l0_idx0(38 downto 38);
-- OL    sum_l0_idx1 <= s_sum_l0_idx1(18 downto 0);
-- OL    c_l0_idx1 <= s_sum_l0_idx1(19 downto 19);
   ----------------Synchro barrier, entering cycle 1----------------
   s_sum_l1_idx1 <=  s_sum_l0_idx1_d1 + c_l0_idx0_d1(0 downto 0);
   sum_l1_idx1 <= s_sum_l1_idx1(18 downto 0);
-- OL    c_l1_idx1 <= s_sum_l1_idx1(19 downto 19);
   R <= sum_l1_idx1(18 downto 0) & sum_l0_idx0_d1(37 downto 0);

   Nc <= s_sum_l0_idx1_d1(18) and s_sum_l0_idx1_d1(17);
end architecture;

--------------------------------------------------------------------------------
--                     FPAdderDualPath_8_47_8_47_8_47400
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPAdderDualPath_8_47_8_47_8_47400 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL     rst : in std_logic;
          X : in  std_logic_vector(8+47+2 downto 0);
          Y : in  std_logic_vector(8+47+2 downto 0);
          R : out  std_logic_vector(8+47+2 downto 0);   
          Nc : out  std_logic);
end entity;

architecture arch of FPAdderDualPath_8_47_8_47_8_47400 is
   component FPAdderDualPath_8_47_8_47_8_47400_DualSubClose is
      port (
-- OL clk : in std_logic;
-- OL        rst : in std_logic;
             X : in  std_logic_vector(49 downto 0);
             Y : in  std_logic_vector(49 downto 0);
             RxMy : out  std_logic_vector(49 downto 0);
             RyMx : out  std_logic_vector(49 downto 0)   );
   end component;

   component FPAdderDualPath_8_47_8_47_8_47400_LZCShifter is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL        rst : in std_logic;
             I : in  std_logic_vector(48 downto 0);
             Count : out  std_logic_vector(5 downto 0);
             O : out  std_logic_vector(48 downto 0)   );
   end component;

   component FPAdderDualPath_8_47_8_47_8_47400_RightShifter is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL        rst : in std_logic;
             X : in  std_logic_vector(47 downto 0);
             S : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(97 downto 0)   );
   end component;

   component FPAdderDualPath_8_47_8_47_8_47400_finalRoundAdd is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL        rst : in std_logic;
             X : in  std_logic_vector(56 downto 0);
             Y : in  std_logic_vector(56 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(56 downto 0);
             Nc : out  std_logic   );
   end component;

   component FPAdderDualPath_8_47_8_47_8_47400_fracAddFar is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL        rst : in std_logic;
             X : in  std_logic_vector(50 downto 0);
             Y : in  std_logic_vector(50 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(50 downto 0);
             Nc : out  std_logic   );
   end component;

signal inX :  std_logic_vector(57 downto 0);
signal inY :  std_logic_vector(57 downto 0);
signal exceptionXSuperiorY : std_logic;
signal exceptionXEqualY : std_logic;
signal signedExponentX :  std_logic_vector(8 downto 0);
signal signedExponentY :  std_logic_vector(8 downto 0);
signal exponentDifferenceXY :  std_logic_vector(8 downto 0);
signal exponentDifferenceYX :  std_logic_vector(7 downto 0);
signal swap : std_logic;
signal newX, newX_d1, newX_d2, newX_d3, newX_d4, newX_d5, newX_d6, newX_d7, newX_d8, newX_d9, newX_d10, newX_d11 :  std_logic_vector(57 downto 0);
signal newY, newY_d1 :  std_logic_vector(57 downto 0);
signal exponentDifference, exponentDifference_d1 :  std_logic_vector(7 downto 0);
signal shiftedOut : std_logic;
signal shiftVal, shiftVal_d1 :  std_logic_vector(5 downto 0);
signal EffSub, EffSub_d1, EffSub_d2, EffSub_d3, EffSub_d4, EffSub_d5, EffSub_d6, EffSub_d7, EffSub_d8, EffSub_d9, EffSub_d10 : std_logic;
signal selectClosePath, selectClosePath_d1, selectClosePath_d2, selectClosePath_d3, selectClosePath_d4, selectClosePath_d5, selectClosePath_d6, selectClosePath_d7, selectClosePath_d8, selectClosePath_d9 : std_logic;
signal sdExnXY, sdExnXY_d1, sdExnXY_d2, sdExnXY_d3, sdExnXY_d4, sdExnXY_d5, sdExnXY_d6, sdExnXY_d7, sdExnXY_d8, sdExnXY_d9, sdExnXY_d10 :  std_logic_vector(3 downto 0);
signal pipeSignY, pipeSignY_d1, pipeSignY_d2, pipeSignY_d3, pipeSignY_d4, pipeSignY_d5, pipeSignY_d6, pipeSignY_d7, pipeSignY_d8, pipeSignY_d9, pipeSignY_d10 : std_logic;
signal fracXClose1 :  std_logic_vector(49 downto 0);
signal fracYClose1 :  std_logic_vector(49 downto 0);
signal fracRClosexMy, fracRClosexMy_d1 :  std_logic_vector(49 downto 0);
signal fracRCloseyMx, fracRCloseyMx_d1 :  std_logic_vector(49 downto 0);
signal fracSignClose, fracSignClose_d1 : std_logic;
signal fracRClose1, fracRClose1_d1 :  std_logic_vector(48 downto 0);
signal resSign, resSign_d1, resSign_d2, resSign_d3, resSign_d4, resSign_d5, resSign_d6, resSign_d7, resSign_d8 : std_logic;
signal nZerosNew, nZerosNew_d1 :  std_logic_vector(5 downto 0);
signal shiftedFrac, shiftedFrac_d1, shiftedFrac_d2 :  std_logic_vector(48 downto 0);
signal roundClose0, roundClose0_d1 : std_logic;
signal resultCloseIsZero0, resultCloseIsZero0_d1 : std_logic;
signal exponentResultClose, exponentResultClose_d1 :  std_logic_vector(9 downto 0);
signal resultBeforeRoundClose :  std_logic_vector(56 downto 0);
signal roundClose : std_logic;
signal resultCloseIsZero : std_logic;
signal fracNewY :  std_logic_vector(47 downto 0);
signal shiftedFracY, shiftedFracY_d1, shiftedFracY_d2 :  std_logic_vector(97 downto 0);
signal sticky, sticky_d1, sticky_d2, sticky_d3 : std_logic;
signal fracYfar :  std_logic_vector(50 downto 0);
signal fracYfarXorOp :  std_logic_vector(50 downto 0);
signal fracXfar :  std_logic_vector(50 downto 0);
signal cInAddFar : std_logic;
signal fracResultfar0, fracResultfar0_d1 :  std_logic_vector(50 downto 0);
signal fracResultFarNormStage :  std_logic_vector(50 downto 0);
signal fracLeadingBits :  std_logic_vector(1 downto 0);
signal fracResultFar1, fracResultFar1_d1 :  std_logic_vector(46 downto 0);
signal fracResultRoundBit : std_logic;
signal fracResultStickyBit : std_logic;
signal roundFar1, roundFar1_d1 : std_logic;
signal expOperationSel :  std_logic_vector(1 downto 0);
signal exponentUpdate :  std_logic_vector(9 downto 0);
signal exponentResultfar0 :  std_logic_vector(9 downto 0);
signal exponentResultFar1, exponentResultFar1_d1 :  std_logic_vector(9 downto 0);
signal resultBeforeRoundFar, resultBeforeRoundFar_d1, resultBeforeRoundFar_d2, resultBeforeRoundFar_d3 :  std_logic_vector(56 downto 0);
signal roundFar, roundFar_d1, roundFar_d2, roundFar_d3 : std_logic;
signal syncClose : std_logic;
signal resultBeforeRound :  std_logic_vector(56 downto 0);
signal round : std_logic;
signal zeroFromClose, zeroFromClose_d1 : std_logic;
signal resultRounded :  std_logic_vector(56 downto 0);
signal syncEffSub : std_logic;
signal syncX :  std_logic_vector(57 downto 0);
signal syncSignY : std_logic;
signal syncResSign : std_logic;
signal UnderflowOverflow :  std_logic_vector(1 downto 0);
signal resultNoExn :  std_logic_vector(57 downto 0);
signal syncExnXY :  std_logic_vector(3 downto 0);
signal exnR :  std_logic_vector(1 downto 0);
signal sgnR : std_logic;
signal expsigR :  std_logic_vector(54 downto 0);

signal NcNewX_a1 : STD_LOGIC ;
signal NcNewX_a2 : STD_LOGIC ;
signal NcNewX_a3 : STD_LOGIC ;
signal NcNewX_a4 : STD_LOGIC ;
signal NcNewX_a5 : STD_LOGIC ;
signal NcPlus    : STD_LOGIC ;
signal NcFinal   : STD_LOGIC ;

begin
   process(clk)
      begin
         if clk'event and clk = '1' then
           if(Enable='1') then
            newX_d1 <=  newX;
            newX_d2 <=  newX_d1;
            newX_d3 <=  newX_d2;
            newX_d4 <=  newX_d3;
            newX_d5 <=  newX_d4;
            newX_d6 <=  newX_d5;
            newX_d7 <=  newX_d6;
            newX_d8 <=  newX_d7;
            newX_d9 <=  newX_d8;
            newX_d10 <=  newX_d9;
            newX_d11 <=  newX_d10;
            newY_d1 <=  newY;
            exponentDifference_d1 <=  exponentDifference;
            shiftVal_d1 <=  shiftVal;
            EffSub_d1 <=  EffSub;
            EffSub_d2 <=  EffSub_d1;
            EffSub_d3 <=  EffSub_d2;
            EffSub_d4 <=  EffSub_d3;
            EffSub_d5 <=  EffSub_d4;
            EffSub_d6 <=  EffSub_d5;
            EffSub_d7 <=  EffSub_d6;
            EffSub_d8 <=  EffSub_d7;
            EffSub_d9 <=  EffSub_d8;
            EffSub_d10 <=  EffSub_d9;
            selectClosePath_d1 <=  selectClosePath;
            selectClosePath_d2 <=  selectClosePath_d1;
            selectClosePath_d3 <=  selectClosePath_d2;
            selectClosePath_d4 <=  selectClosePath_d3;
            selectClosePath_d5 <=  selectClosePath_d4;
            selectClosePath_d6 <=  selectClosePath_d5;
            selectClosePath_d7 <=  selectClosePath_d6;
            selectClosePath_d8 <=  selectClosePath_d7;
            selectClosePath_d9 <=  selectClosePath_d8;
            sdExnXY_d1 <=  sdExnXY;
            sdExnXY_d2 <=  sdExnXY_d1;
            sdExnXY_d3 <=  sdExnXY_d2;
            sdExnXY_d4 <=  sdExnXY_d3;
            sdExnXY_d5 <=  sdExnXY_d4;
            sdExnXY_d6 <=  sdExnXY_d5;
            sdExnXY_d7 <=  sdExnXY_d6;
            sdExnXY_d8 <=  sdExnXY_d7;
            sdExnXY_d9 <=  sdExnXY_d8;
            sdExnXY_d10 <=  sdExnXY_d9;
            pipeSignY_d1 <=  pipeSignY;
            pipeSignY_d2 <=  pipeSignY_d1;
            pipeSignY_d3 <=  pipeSignY_d2;
            pipeSignY_d4 <=  pipeSignY_d3;
            pipeSignY_d5 <=  pipeSignY_d4;
            pipeSignY_d6 <=  pipeSignY_d5;
            pipeSignY_d7 <=  pipeSignY_d6;
            pipeSignY_d8 <=  pipeSignY_d7;
            pipeSignY_d9 <=  pipeSignY_d8;
            pipeSignY_d10 <=  pipeSignY_d9;
            fracRClosexMy_d1 <=  fracRClosexMy;
            fracRCloseyMx_d1 <=  fracRCloseyMx;
            fracSignClose_d1 <=  fracSignClose;
            fracRClose1_d1 <=  fracRClose1;
            resSign_d1 <=  resSign;
            resSign_d2 <=  resSign_d1;
            resSign_d3 <=  resSign_d2;
            resSign_d4 <=  resSign_d3;
            resSign_d5 <=  resSign_d4;
            resSign_d6 <=  resSign_d5;
            resSign_d7 <=  resSign_d6;
            resSign_d8 <=  resSign_d7;
            nZerosNew_d1 <=  nZerosNew;
            shiftedFrac_d1 <=  shiftedFrac;
            shiftedFrac_d2 <=  shiftedFrac_d1;
            roundClose0_d1 <=  roundClose0;
            resultCloseIsZero0_d1 <=  resultCloseIsZero0;
            exponentResultClose_d1 <=  exponentResultClose;
            shiftedFracY_d1 <=  shiftedFracY;
            shiftedFracY_d2 <=  shiftedFracY_d1;
            sticky_d1 <=  sticky;
            sticky_d2 <=  sticky_d1;
            sticky_d3 <=  sticky_d2;
            fracResultfar0_d1 <=  fracResultfar0;
            fracResultFar1_d1 <=  fracResultFar1;
            roundFar1_d1 <=  roundFar1;
            exponentResultFar1_d1 <=  exponentResultFar1;
            resultBeforeRoundFar_d1 <=  resultBeforeRoundFar;
            resultBeforeRoundFar_d2 <=  resultBeforeRoundFar_d1;
            resultBeforeRoundFar_d3 <=  resultBeforeRoundFar_d2;
            roundFar_d1 <=  roundFar;
            roundFar_d2 <=  roundFar_d1;
            roundFar_d3 <=  roundFar_d2;
            zeroFromClose_d1 <=  zeroFromClose;
           end if;
         end if;
      end process;
-- Exponent difference and swap  --
   inX <= X;
   inY <= Y;
   exceptionXSuperiorY <= '1' when inX(57 downto 56) >= inY(57 downto 56) else '0';
   exceptionXEqualY <= '1' when inX(57 downto 56) = inY(57 downto 56) else '0';
   signedExponentX <= "0" & inX(54 downto 47);
   signedExponentY <= "0" & inY(54 downto 47);
   exponentDifferenceXY <= signedExponentX - signedExponentY ;
   exponentDifferenceYX <= signedExponentY(7 downto 0) - signedExponentX(7 downto 0);
   swap <= (exceptionXEqualY and exponentDifferenceXY(8)) or (not(exceptionXSuperiorY));
   newX <= inY when swap = '1' else inX;
   newY <= inX when swap = '1' else inY;
   exponentDifference <= exponentDifferenceYX when swap = '1' else exponentDifferenceXY(7 downto 0);
   shiftedOut <= exponentDifference(7) or exponentDifference(6);
   shiftVal <= exponentDifference(5 downto 0) when shiftedOut='0'
          else CONV_STD_LOGIC_VECTOR(50,6) ;
   ----------------Synchro barrier, entering cycle 1----------------
   EffSub <= newX_d1(55) xor newY_d1(55);
   selectClosePath <= EffSub when exponentDifference_d1(7 downto 1) = (7 downto 1 => '0') else '0';
   sdExnXY <= newX_d1(57 downto 56) & newY_d1(57 downto 56);
   pipeSignY <= newY_d1(55);

-- Close Path --
   fracXClose1 <= "01" & newX_d1(46 downto 0) & '0';
   with exponentDifference_d1(0) select
   fracYClose1 <=  "01" & newY_d1(46 downto 0) & '0' when '0',
                  "001" & newY_d1(46 downto 0)       when others;
   DualSubO: FPAdderDualPath_8_47_8_47_8_47400_DualSubClose  -- pipelineDepth=0 maxInDelay=0
      port map (
-- OL clk  => clk,
-- OL                 rst  => rst,
                 RxMy => fracRClosexMy,
                 RyMx => fracRCloseyMx,
                 X => fracXClose1,
                 Y => fracYClose1);
   ----------------Synchro barrier, entering cycle 2----------------
   fracSignClose <= fracRClosexMy_d1(49);
   fracRClose1 <= fracRClosexMy_d1(48 downto 0) when fracSignClose='0' else fracRCloseyMx_d1(48 downto 0);
   ----------------Synchro barrier, entering cycle 3----------------
   resSign <= '0' when selectClosePath_d2='1' and fracRClose1_d1 = (48 downto 0 => '0') else
             newX_d3(55) xor (selectClosePath_d2 and fracSignClose_d1);
   LZC_component: FPAdderDualPath_8_47_8_47_8_47400_LZCShifter  -- pipelineDepth=5 maxInDelay=0
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 Count => nZerosNew,
                 I => fracRClose1_d1,
                 O => shiftedFrac);
   ----------------Synchro barrier, entering cycle 8----------------
   ----------------Synchro barrier, entering cycle 9----------------
   roundClose0 <= shiftedFrac_d1(0) and shiftedFrac_d1(1);
   resultCloseIsZero0 <= '1' when nZerosNew_d1 = CONV_STD_LOGIC_VECTOR(49, 6) else '0';
   exponentResultClose <= ("00" & newX_d9(54 downto 47)) - (CONV_STD_LOGIC_VECTOR(0,4) & nZerosNew_d1);
   ----------------Synchro barrier, entering cycle 10----------------
   resultBeforeRoundClose <= exponentResultClose_d1(9 downto 0) & shiftedFrac_d2(47 downto 1);
   roundClose <= roundClose0_d1;
   resultCloseIsZero <= resultCloseIsZero0_d1;

-- Far Path --
   ---------------- cycle 1----------------
   fracNewY <= '1' & newY_d1(46 downto 0);
   RightShifterComponent: FPAdderDualPath_8_47_8_47_8_47400_RightShifter  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                  rst  => rst,
                 R => shiftedFracY,
                 S => shiftVal_d1,
                 X => fracNewY);
   ----------------Synchro barrier, entering cycle 3----------------
   sticky <= '0' when (shiftedFracY_d1(47 downto 0)=CONV_STD_LOGIC_VECTOR(0,47)) else '1';
   ----------------Synchro barrier, entering cycle 4----------------
   fracYfar <= "0" & shiftedFracY_d2(97 downto 48);
   fracYfarXorOp <= fracYfar xor (50 downto 0 => EffSub_d3);
   fracXfar <= "01" & (newX_d4(46 downto 0)) & "00";
   cInAddFar <= EffSub_d3 and not sticky_d1;
   fracAdderFar: FPAdderDualPath_8_47_8_47_8_47400_fracAddFar  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                  rst  => rst,
                 Cin => cInAddFar,
                 R => fracResultfar0,
                 X => fracXfar,
                 Y => fracYfarXorOp,
                 Nc => NcPlus);
   ----------------Synchro barrier, entering cycle 5----------------
   ----------------Synchro barrier, entering cycle 6----------------
   -- 2-bit normalisation
   fracResultFarNormStage <= fracResultfar0_d1;
   fracLeadingBits <= fracResultFarNormStage(50 downto 49) ;
   fracResultFar1 <=
           fracResultFarNormStage(47 downto 1)  when fracLeadingBits = "00"
      else fracResultFarNormStage(48 downto 2)  when fracLeadingBits = "01"
      else fracResultFarNormStage(49 downto 3);
   fracResultRoundBit <=
           fracResultFarNormStage(0)     when fracLeadingBits = "00"
      else fracResultFarNormStage(1)    when fracLeadingBits = "01"
      else fracResultFarNormStage(2) ;
   fracResultStickyBit <=
           sticky_d3     when fracLeadingBits = "00"
      else fracResultFarNormStage(0) or  sticky_d3   when fracLeadingBits = "01"
      else fracResultFarNormStage(1) or fracResultFarNormStage(0) or sticky_d3;
   roundFar1 <= fracResultRoundBit and (fracResultStickyBit or fracResultFar1(0));
   expOperationSel <= "11" when fracLeadingBits = "00" -- add -1 to exponent
               else   "00" when fracLeadingBits = "01" -- add 0 
               else   "01";                              -- add 1
   exponentUpdate <= (9 downto 1 => expOperationSel(1)) & expOperationSel(0);
   exponentResultfar0<="00" & (newX_d6(54 downto 47));
   exponentResultFar1 <= exponentResultfar0 + exponentUpdate;
   ----------------Synchro barrier, entering cycle 7----------------
   resultBeforeRoundFar <= exponentResultFar1_d1 & fracResultFar1_d1;
   roundFar <= roundFar1_d1;

-- Synchronization of both paths --
   ---------------- cycle 7----------------
   ----------------Synchro barrier, entering cycle 10----------------
   syncClose <= selectClosePath_d9;
   with syncClose select
   resultBeforeRound <= resultBeforeRoundClose when '1',
                        resultBeforeRoundFar_d3   when others;
   with syncClose select
   round <= roundClose when '1',
            roundFar_d3   when others;
   zeroFromClose <= syncClose and resultCloseIsZero;

-- Rounding --
   finalRoundAdder: FPAdderDualPath_8_47_8_47_8_47400_finalRoundAdd  -- pipelineDepth=1 maxInDelay=9.4872e-10
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 Cin => round,
                 R => resultRounded,
                 X => resultBeforeRound,
                 Y => (56 downto 0 => '0'), 
                 Nc => NcFinal );
   syncEffSub <= EffSub_d10;
   syncX <= newX_d11;
   syncSignY <= pipeSignY_d10;
   syncResSign <= resSign_d8;
   UnderflowOverflow <= resultRounded(56 downto 55);
   with UnderflowOverflow select
   resultNoExn(57 downto 56) <=   (not zeroFromClose_d1) & "0" when "01", -- overflow
                                 "00" when "10" | "11",  -- underflow
                                 "0" &  not zeroFromClose_d1  when others; -- normal 
   resultNoExn(55 downto 0) <= syncResSign & resultRounded(54 downto 0);
   syncExnXY <= sdExnXY_d10;
   -- Exception bits of the result
   with syncExnXY select -- remember that ExnX > ExnY 
      exnR <= resultNoExn(57 downto 56) when "0101",
              "1" & syncEffSub          when "1010",
              "11"                      when "1110",
              syncExnXY(3 downto 2)     when others;
   -- Sign bit of the result
   with syncExnXY select
      sgnR <= resultNoExn(55)         when "0101",
              syncX(55) and syncSignY when "0000",
              syncX(55)               when others;
   -- Exponent and significand of the result
   with syncExnXY select
      expsigR <= resultNoExn(54 downto 0)   when "0101" ,
                 syncX(54 downto  0)        when others; -- 0100, or at least one NaN or one infty 
   R <= exnR & sgnR & expsigR;

NcNewX_a1 <= newX_d2(56) and newX_d2(57)and newX_d3(56) and newX_d3(57) and newX_d4(56) and newX_d4(57);
NcNewX_a2 <= newX_d5(56) and newX_d5(57)and newX_d6(56) and newX_d6(57) and newX_d7(56) and newX_d7(57);
NcNewX_a3 <= newX_d8(56) and newX_d8(57)and newX_d9(56) and newX_d9(57) and newX_d10(56) and newX_d10(57);
NcNewX_a4 <= newX_d11(56) and newX_d11(57) and shiftedFrac_d1(48) and NcPlus;
NcNewX_a5 <= EffSub_d4 and EffSub_d5 and EffSub_d6 and EffSub_d7 and EffSub_d8 and EffSub_d9 and EffSub_d10;

Nc <= NcNewX_a1 and NcNewX_a2 and NcNewX_a3 and NcNewX_a4 and NcNewX_a5 and NcFinal;


end architecture;

