
library IEEE;
use IEEE.std_logic_1164.all;

package TransCtrlPack is

  constant FlitWidth : natural :=16;
  
end TransCtrlPack;
