--------------------------------------------------------------------------------
--                             firstExpTable_9_52
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity firstExpTable_9_52 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(51 downto 0)   );
end entity;

architecture arch of firstExpTable_9_52 is
   -- Build a 2-D array type for the RoM
   subtype word_t is std_logic_vector(51 downto 0);
   type memory_t is array(0 to 511) of word_t;
   function init_rom
      return memory_t is 
      variable tmp : memory_t := (
   "1000000000000000000000000000000000000000000000000000",
   "1000000001000000000100000000001010101011000000000001",
   "1000000010000000010000000001010101011010101010111100",
   "1000000011000000100100000100100000011011000010000010",
   "1000000100000001000000001010101100000000001000100011",
   "1000000101000001100100010100111000100110000100110000",
   "1000000110000010010000100100000110110001000000111011",
   "1000000111000011000100111001010111001101001100011000",
   "1000001000000100000001010101101010101110111100011101",
   "1000001001000101000101111010000010010010101101100001",
   "1000001010000110010010100111011110111101000100000011",
   "1000001011000111100111011111000001111010101101100101",
   "1000001100001001000100100001101100100000100001101111",
   "1000001101001010101001110000100000001011100011010000",
   "1000001110001100010111001100011110100001000001000010",
   "1000001111001110001100110110101001001110010111001010",
   "1000010000010000001010110000000010001001001111110110",
   "1000010001010010010000111001101011001111100100100110",
   "1000010010010100011111010100100110100111011111001000",
   "1000010011010110110110000001110110011111011010011101",
   "1000010100011001010101000010011101001110000011111011",
   "1000010101011011111100010111011101010010011100001101",
   "1000010110011110101100000001111001010011111000011001",
   "1000010111100001100100000010110100000010000011000001",
   "1000011000100100100100011011010000010100111101000110",
   "1000011001100111101101001100010001001100111111001000",
   "1000011010101010111110010110111001110010111010001111",
   "1000011011101110010111111100001101010111111001001001",
   "1000011100110001111001111101001111010101100001001111",
   "1000011101110101100100011011000011001101110011101000",
   "1000011110111001010111010110101100101011001110001110",
   "1000011111111101010010110001001111100000101100110000",
   "1000100001000001010110101011101111101001101001110111",
   "1000100010000101100011000111010001001010000000001000",
   "1000100011001001111000000100111000001110001011001011",
   "1000100100001110010101100101101001001011001000101100",
   "1000100101010010111011101010101000011110011001100010",
   "1000100110010111101010010100111010101110000010110011",
   "1000100111011100100001100101100100101000101110110101",
   "1000101000100001100001011101101011000101101110011001",
   "1000101001100110101001111110010011000100111001101011",
   "1000101010101011111011001000100001101110110001011001",
   "1000101011110001010100111101011100010100011111110110",
   "1000101100110110110111011110001000001111111010000100",
   "1000101101111100100010101011101011000011100000110101",
   "1000101111000010010110100111001010011010100001110000",
   "1000110000001000010011010001101100001000111000011010",
   "1000110001001110011000101100010110001011001111011101",
   "1000110010010100100110111000001110100111000001100111",
   "1000110011011010111101110110011011101010011010110110",
   "1000110100100001011101101000000011101100011001011110",
   "1000110101101000000110001110001101001100101111001101",
   "1000110110101110110111101001111110110100000010010001",
   "1000110111110101110001111100011111010011101110100011",
   "1000111000111100110101000110110101100110000110101000",
   "1000111010000100000001001010001000101110010100111110",
   "1000111011001011010110000111011111111000011100111101",
   "1000111100010010110100000000000010011001011100000001",
   "1000111101011010011010110100110111101111001010110101",
   "1000111110100010001010100111000111100000011110010010",
   "1000111111101010000011010111111001011101001000101111",
   "1001000000110010000101001000010101011101111011000100",
   "1001000001111010001111111001100011100100100101110010",
   "1001000011000010100011101100101011111011111010001110",
   "1001000100001011000000100010110110110111101011100110",
   "1001000101010011100110011101001100110100110000001100",
   "1001000110011100010101011100110110011001000010011010",
   "1001000111100101001101100010111100010011100010000010",
   "1001001000101110001110110000100111011100010101001101",
   "1001001001110111011001000111000000110100101001101111",
   "1001001011000000101100100111010001100110110110000111",
   "1001001100001010001001010010100011000110011010101010",
   "1001001101010011101111001001111110110000000010110010",
   "1001001110011101011110001110101110001001100101111111",
   "1001001111100111010110100001111011000010001001001000",
   "1001010000110001011000000100101111010001111111011111",
   "1001010001111011100010111000010100111010101011111111",
   "1001010011000101110110111101110110000111000010010011",
   "1001010100010000010100010110011101001011001000000011",
   "1001010101011010111011000011010100100100010101111100",
   "1001010110100101101011000101100110111001011000111101",
   "1001010111110000100100011110011110111010010011011100",
   "1001011000111011100111001111000111100000011110011001",
   "1001011010000110110011011000101011101110101010100011",
   "1001011011010010001000111100010110110001000001100100",
   "1001011100011101100111111011010011111101000111001101",
   "1001011101101001010000010110101110110001111010100001",
   "1001011110110101000010001111110010110111110111000011",
   "1001100000000000111101100111101100000000110101111100",
   "1001100001001101000010011111100110001000001111001011",
   "1001100010011001010000111000101101010010111010110010",
   "1001100011100101101000110100001101101111010001111101",
   "1001100100110010001010010011010011110101010000010100",
   "1001100101111110110101010111001100000110010101000100",
   "1001100111001011101010000001000011001101100100001001",
   "1001101000011000101000010010000101111111100111100011",
   "1001101001100101110000001011100001011010110000011011",
   "1001101010110011000001101110100010100110111000010001",
   "1001101100000000011100111100010110110101100010001111",
   "1001101101001110000001110110001011100001111100001110",
   "1001101110011011110000011101001110010001000000001001",
   "1001101111101001101000110010101100110001010101001011",
   "1001110000110111101010110111110100111011010000110111",
   "1001110010000101110110101101110100110000111000011101",
   "1001110011010100001100010101111010011110000010000011",
   "1001110100100010101011110001010100011000010101110101",
   "1001110101110001010101000001010000111111001111010100",
   "1001110111000000001000000110111110111011111110100010",
   "1001111000001111000101000011101101000001101001010101",
   "1001111001011110001011111000101010001101001100100001",
   "1001111010101101011100100111000101100101011101001001",
   "1001111011111100110111010000001110011011001001110001",
   "1001111101001100011011110101010100001000111011100110",
   "1001111110011100001010010111100110010011010111110110",
   "1001111111101100000010111000010100101001000000111001",
   "1010000000111100000101011000101111000010010111100100",
   "1010000010001100010001111010000101100001111100011001",
   "1010000011011100101000011101101000010100010000110100",
   "1010000100101101001001000100100111101111111000100000",
   "1010000101111101110011110000010100010101011010100001",
   "1010000111001110101000100001111110101111100010101100",
   "1010001000011111100111011010110111110011000010110010",
   "1010001001110000110000011100010000011110110011110010",
   "1010001011000010000011100111011001111011110111001100",
   "1010001100010011100000111101100101011101011000010000",
   "1010001101100101001000100000000100100000101101010001",
   "1010001110110110111010010000001000101101011000110100",
   "1010010000001000110110001111000011110101001011000100",
   "1010010001011010111100011110000111110100000011000011",
   "1010010010101101001100111110100110110000001111111101",
   "1010010011111111100111110001110010111010010010010110",
   "1010010101010010001100111000111110101100111101100010",
   "1010010110100100111100010101011100101101011000110100",
   "1010010111110111110110001000011111101011000000110000",
   "1010011001001010111010010011011010011111101000100000",
   "1010011010011110001000110111100000001111011011000111",
   "1010011011110001100001110110000100001000111100110000",
   "1010011101000101000101010000011001100101001100000111",
   "1010011110011000110011000111110100000111100011101000",
   "1010011111101100101011011101100111011101111010110100",
   "1010100001000000101110010011000111100000100111100110",
   "1010100010010100111011101001101000010010011111100110",
   "1010100011101001010011100010011110000000111001011010",
   "1010100100111101110101111110111101000011101101111111",
   "1010100110010010100011000000011001111101011001111100",
   "1010100111100111011010101000001001011010111110110100",
   "1010101000111100011100110111100000010100000100011111",
   "1010101010010001101001101111110011101010111010011001",
   "1010101011100111000001010010011000101100011000111110",
   "1010101100111100100011100000100100110000000010111001",
   "1010101110010010010000011011101101011000000110011111",
   "1010101111101000001000000101001000010001011110111110",
   "1010110000111110001010011110001011010011110101111000",
   "1010110010010100010111101000001100100001100100011000",
   "1010110011101010101111100100100010000111110100100111",
   "1010110101000001010010010100100010011110100011000001",
   "1010110110010111111111111001100100001000011111101101",
   "1010110111101110111000010100111101110011001111110100",
   "1010111001000101111011101000000110010111001110111000",
   "1010111010011101001001110100010100110111110000001000",
   "1010111011110100100010111011000000100010111111111011",
   "1010111101001100000110111101100000110010000101000010",
   "1010111110100011110101111101001101001001000010000101",
   "1010111111111011101111111011011101010110110110111001",
   "1011000001010011110100111001101001010101100001110100",
   "1011000010101100000100111001001001001010000001001011",
   "1011000100000100011111111011010101000100010100100011",
   "1011000101011101000110000001100101011111011110010001",
   "1011000110110101110111001101010011000001100100101100",
   "1011001000001110110011011111110110011011110011101010",
   "1011001001100111111010111010101000101010011101110100",
   "1011001011000001001101011111000010110100111110000101",
   "1011001100011010101011001110011110001101111000111110",
   "1011001101110100010100001010010100010010111110000011",
   "1011001111001110001000010011111110101101001001010000",
   "1011010000101000000111101100110111010000100100010111",
   "1011010010000010010010010110010111111100101000011001",
   "1011010011011100101000010001111010111011111110111110",
   "1011010100110111001001100000111010100100100011110001",
   "1011010110010001110110000100110001010111100101111000",
   "1011010111101100101101111110111010000001101001010001",
   "1011011001000111110001010000101111011010101000001110",
   "1011011010100010111111111011101100100101110100101011",
   "1011011011111110011010000001001100110001111001101101",
   "1011011101011001111111100010101011011000111100111011",
   "1011011110110101110000100001100100000000011111111100",
   "1011100000010001101100111111010010011001100001110000",
   "1011100001101101110100111101010010100000100000001110",
   "1011100011001010001000011101000000011101011001011101",
   "1011100100100110100111011111111000100011101101010010",
   "1011100110000011010010000111010111010010011110101101",
   "1011100111100000001000010100111001010100010101010110",
   "1011101000111101001010001001111011011111011110110101",
   "1011101010011010010111100111111010110101110000010101",
   "1011101011110111110000110000010100100100100111111100",
   "1011101101010101010101100100100110000101001110001101",
   "1011101110110011000110000110001100111100010111100000",
   "1011110000010001000010010110100110111010100101100101",
   "1011110001101111001010010111010001111100001000111100",
   "1011110011001101011110001001101100001001000010011010",
   "1011110100101011111101101111010011110101000100011111",
   "1011110110001010101001001001100111011111110100111100",
   "1011110111101001100000011010000101110100101110001011",
   "1011111001001000100011100010001101101011000000110101",
   "1011111010100111110010100011011110000101110101000111",
   "1011111100000111001101011111010110010100001100011010",
   "1011111101100110110100010111010101110001000010101111",
   "1011111111000110100111001100111100000011010000001110",
   "1100000000100110100110000001101000111101101010100011",
   "1100000010000110110000110110111100011111000110100100",
   "1100000011100111000111101110010110110010011001101110",
   "1100000101000111101010101001011000001110011011100001",
   "1100000110101000011001101001100001010110000111001000",
   "1100001000001001010100110000010010111000011100110100",
   "1100001001101010011011111111001101110000100011011101",
   "1100001011001011101111010111110011000101101010001001",
   "1100001100101101001110111011100100001011001001100011",
   "1100001110001110111010101100000010100000100101100101",
   "1100001111110000110010101010101111110001101110110101",
   "1100010001010010110110111001001101110110100100001001",
   "1100010010110101000111011000111110110011010100000111",
   "1100010100010111100100001011100100111000011110101001",
   "1100010101111010001101010010100010100010110110011100",
   "1100010111011101000010101111011010011011100010100110",
   "1100011001000000000100100011101111011000000000001000",
   "1100011010100011010010110001000100011010000011011111",
   "1100011100000110101101011000111100101111111010000111",
   "1100011101101010010100011100111011110100001100000010",
   "1100011111001110000111111110100101001101111101011000",
   "1100100000110010000111111111011100110000101111111001",
   "1100100010010110010100100001000110011100100100100101",
   "1100100011111010101101100101000110011101111101010000",
   "1100100101011111010011001101000001001101111110000000",
   "1100100111000100000101011010011011010010001110111001",
   "1100101000101001000100001110111001011100111101011110",
   "1100101010001110001111101100000000101100111110010110",
   "1100101011110011100111110011010110001101101110101111",
   "1100101101011001001100100110011111010111010110001000",
   "1100101110111110111110000111000001101110100111110010",
   "1100110000100100111100010110100011000101000100011001",
   "1100110010001011000111010110101001011000111011100110",
   "1100110011110001011111001000111010110101001101101000",
   "1100110101011000000011101110111101110001101100111001",
   "1100110110111110110101001010011000110010111111100100",
   "1100111000100101110011011100110010101010100001001110",
   "1100111010001100111110100111110010010110100100010111",
   "1100111011110100010110101100111111000010010100001010",
   "1100111101011011111011101110000000000101110101111011",
   "1100111111000011101101101100011101000110001010110011",
   "1101000000101011101100101001111101110101010001011001",
   "1101000010010011111000101000001010010010000111010110",
   "1101000011111100010001101000101010101000101010111110",
   "1101000101100100110111101101000111010001111100111100",
   "1101000111001101101010110111001000110100000001110100",
   "1101001000110110101011001000011000000010000011110000",
   "1101001010011111111000100010011101111100010100001001",
   "0100110110100010110010111111000110111110010110000010",
   "0100110111001001101001110000110110101110111110000100",
   "0100110111110000100101011001110000001001110000110111",
   "0100111000010111100101111010011010001010010111011010",
   "0100111000111110101011010011011011110001010010011000",
   "0100111001100101110101100101011100000011111010111000",
   "0100111010001101000100110001000010001100100010111100",
   "0100111010110100011000110110110101011010010110001110",
   "0100111011011011110001110111011101000001011010100100",
   "0100111100000011001111110011100000011010110000101010",
   "0100111100101010110010101011100111000100010100100110",
   "0100111101010010011010100000011000100000111110100010",
   "0100111101111010000111010010011100011000100011010010",
   "0100111110100001111001000010011010010111110100111111",
   "0100111111001001101111110000111010010000100011101000",
   "0100111111110001101011011110100011111001011101110010",
   "0101000000011001101100001011111111001110010001001010",
   "0101000001000001110001111001110100001111101011001101",
   "0101000001101001111100101000101011000011011001110101",
   "0101000010010010001100011001001011110100001011111011",
   "0101000010111010100001001011111110110001110010000100",
   "0101000011100010111011000001101100010000111111000110",
   "0101000100001011011001111010111100101011101000110010",
   "0101000100110011111101111000011000100000101000011100",
   "0101000101011100100110111010101000010011111011100010",
   "0101000110000101010101000010010100101110100100011000",
   "0101000110101110001000010000000110011110101010101111",
   "0101000111010111000000100100100110010111011100011010",
   "0101000111111111111110000000011101010001001101111101",
   "0101001000101001000000100100010100001001011011010011",
   "0101001001010010001000010000110100000010101000010110",
   "0101001001111011010101000110100110000100100001101001",
   "0101001010100100100111000110010011011011111101000010",
   "0101001011001101111110010000100101011010111010010010",
   "0101001011110111011010100110000101011000100011101101",
   "0101001100100000111100000111011100110001001110110111",
   "0101001101001010100010110101010101000110011101001100",
   "0101001101110100001110110000010111111110111100100111",
   "0101001110011101111111111001001111000110101000001110",
   "0101001111000111110110010000100100001110101000111100",
   "0101001111110001110001110111000001001101010110001010",
   "0101010000011011110010101101001111111110010110010111",
   "0101010001000101111000110011111010100010011111110111",
   "0101010001110000000100001011101010111111111001010111",
   "0101010010011010010100110101001011100001111010101100",
   "0101010011000100101010110001000110011001001101011001",
   "0101010011101111000110000000000101111011101101011101",
   "0101010100011001100110100010110100100100101001111010",
   "0101010101000100001100011001111100110100100101100100",
   "0101010101101110110111100110001001010001010111100110",
   "0101010110011001101000001000000100100110001100001111",
   "0101010111000100011110000000011001100011100101011111",
   "0101010111101111011001001111110010111111011011101110",
   "0101011000011010011001110110111011110100111110011010",
   "0101011001000101011111110110011111000100110100101110",
   "0101011001110000101011001111000111110100111110010010",
   "0101011010011011111100000001100001010000110011110010",
   "0101011011000111010010001110010110101001000111101011",
   "0101011011110010101101110110010011010100000110110101",
   "0101011100011110001110111010000010101101011001010010",
   "0101011101001001110101011010010000010110000010110100",
   "0101011101110101100001010111100111110100100011101101",
   "0101011110100001010010110010110100110100111001010111",
   "0101011111001101001001101100100011001000011111000011",
   "0101011111111001000110000101011110100110001110100100",
   "0101100000100101000111111110010011001010100000111000",
   "0101100001010001001111010111101100110111001110110111",
   "0101100001111101011100010010010111110011110010000000",
   "0101100010101001101110101111000000001101000101000000",
   "0101100011010110000110101110010010010101100100100100",
   "0101100100000010100100010000111010100101010000000001",
   "0101100100101111000111010111100101011001101010000100",
   "0101100101011011110000000010111111010101111001011011",
   "0101100110001000011110010011110101000010101001100011",
   "0101100110110101010010001010110011001110001011010111",
   "0101100111100010001011101000100110101100010101110111",
   "0101101000001111001010101101111100010110100110111100",
   "0101101000111100001111011011100001001100000011111110",
   "0101101001101001011001110010000010010001011010100111",
   "0101101010010110101001110010001100110001000001011010",
   "0101101011000011111111011100101101111010111000100111",
   "0101101011110001011010110010010011000100101010110010",
   "0101101100011110111011110011101001101001101101100101",
   "0101101101001100100010100001011111001011000010011001",
   "0101101101111010001110111100100001001111010111001000",
   "0101101110101000000001000101011101100011000110110111",
   "0101101111010101111000111101000001111000011010101000",
   "0101110000000011110110100011111100000111001010000001",
   "0101110000110001111001111010111010001100111100000010",
   "0101110001100000000011000010101010001101000111101011",
   "0101110010001110010001111011111010010000110100110010",
   "0101110010111100100110100111011000100110111100101001",
   "0101110011101011000001000101110011100100001010110011",
   "0101110100011001100001010111111001100010111101101111",
   "0101110101001000000111011110011001000011100111100111",
   "0101110101110110110011011010000000101100001110111110",
   "0101110110100101100101001011011111001000101111100000",
   "0101110111010100011100110011100011001010111010101110",
   "0101111000000011011010010010111011101010011000110001",
   "0101111000110010011101101010010111100100101001000110",
   "0101111001100001100110111010100101111101000011001011",
   "0101111010010000110110000100010101111100110111010100",
   "0101111011000000001011001000010110110011001111010101",
   "0101111011101111100110000111010111110101001111010001",
   "0101111100011111000111000010001000011101110110001111",
   "0101111101001110101101111001011000001101111111000010",
   "0101111101111110011010101101110110101100100000111111",
   "0101111110101110001101100000010011100110010000101000",
   "0101111111011110000110010001011110101110000000011110",
   "0110000000001110000101000010000111111100100001101111",
   "0110000000111110001001110010111111010000100101001010",
   "0110000001101110010100100100110100101110111011101001",
   "0110000010011110100101011000011000100010010111000101",
   "0110000011001110111100001110011010111011101011001000",
   "0110000011111111011001000111101100010001101101110111",
   "0110000100101111111100000100111101000001011000100111",
   "0110000101100000100101000110111101101101101000101110",
   "0110000110010001010100001110011110111111100000010000",
   "0110000111000010001001011100010001100110000110110010",
   "0110000111110011000100110001000110010110101010001100",
   "0110001000100100000110001101101110001100011111010101",
   "0110001001010101001101110010111010001001000010111010",
   "0110001010000110011011100001011011010011111010001011",
   "0110001010110111101111011010000010111010110011101110",
   "0110001011101001001001011101100010010001101000001101",
   "0110001100011010101001101100101010110010011011001100",
   "0110001101001100010000001000001101111101011011111001",
   "0110001101111101111100110000111101011001000101111010",
   "0110001110101111101111100111101010110010000010000011",
   "0110001111100001101000101101000111111011000111000101",
   "0110010000010011101000000010000110101101011010100010",
   "0110010001000101101101100111011001001000010001011100",
   "0110010001110111111001011101110001010001010001001011",
   "0110010010101010001011100110000001010100010000001011",
   "0110010011011100100100000000111011100011010110101111",
   "0110010100001111000010101111010010010110111111110111",
   "0110010101000001100111110001111000001101111001111101",
   "0110010101110100010011001001011111101101000111101011",
   "0110010110100111000100110110111011100000000000101101",
   "0110010111011001111100111010111110011000010010100011",
   "0110011000001100111011010110011011001110000001010101",
   "0110011001000000000000001010000100111111101000100011",
   "0110011001110011001011010110101110110001111011111011",
   "0110011010100110011100111101001011110000001000001100",
   "0110011011011001110100111110001111001011110011110110",
   "0110011100001101010011011010101100011101000000000001",
   "0110011101000000111000010011010111000010001001010000",
   "0110011101110100100011101001000010100000001000010000",
   "0110011110101000010101011100100010100010010010110010",
   "0110011111011100001101101110101010111010011100011010",
   "0110100000010000001100100000001111100000110111010100",
   "0110100001000100010001110010000100010100010101001010",
   "0110100001111000011101100100111101011010000111110100",
   "0110100010101100101111111001101110111110000010010001",
   "0110100011100001001000110001001101010010011001010101",
   "0110100100010101101000001100001100110000000100100101",
   "0110100101001010001110001011100001110110011111000010",
   "0110100101111110111010110000000001001011101000001000",
   "0110100110110011101101111010011111011100000100011010",
   "0110100111101000100111101011110001011010111110011010",
   "0110101000011101101000000100101100000010000111011111",
   "0110101001010010101111000110000100010001111000101000",
   "0110101010000111111100110000101111010001010011010001",
   "0110101010111101010001000101100010001110000010001010",
   "0110101011110010101100000101010010011100011010001011",
   "0110101100101000001101110000110101010111011011000111",
   "0110101101011101110110001001000000100000110000100111",
   "0110101110010011100101001110101001100000110010111010",
   "0110101111001001011011000010100110000110100111101101",
   "0110101111111111010111100101101100001000000011000010",
   "0110110000110101011010111000110001100001101000000011",
   "0110110001101011100100111100101100010110101001111010",
   "0110110010100001110101110010010010110001001100100110",
   "0110110011011000001101011010011011000010000101110011",
   "0110110100001110101011110101111011100000111101101100",
   "0110110101000101010001000101101010101100001111111000",
   "0110110101111011111101001010011111001001001100001010",
   "0110110110110010110000000101001111100011110111011010",
   "0110110111101001101001110110110010101111001100011110",
   "0110111000100000101010011111111111100100111100111101",
   "0110111001010111110010000001101101000101110010001010",
   "0110111010001111000000011100110010011001001101110110",
   "0110111011000110010101110010000110101101101011001010",
   "0110111011111101110010000010100001011000011111100001",
   "0110111100110101010101001110111001110101111011011001",
   "0110111101101100111111011000000111101001001011001111",
   "0110111110100100110000011111000010011100011000010101",
   "0110111111011100101000100100100010000000101001101100",
   "0111000000010100100111101001011110001110000100110111",
   "0111000001001100101101101110101111000011101110111000",
   "0111000010000100111010110101001100100111101101000011",
   "0111000010111101001110111101101111000111000101111100",
   "0111000011110101101010001001001110110110000010001000",
   "0111000100101110001100011000100100001111101101001110",
   "0111000101100110110101101100100111110110010110100110",
   "0111000110011111100110000110010010010011010010011001",
   "0111000111011000011101100110011100010110111010010110",
   "0111001000010001011100001101111110111000101110101101",
   "0111001001001010100001111101110010110111010111000011",
   "0111001010000011101110110110110001011000100011010011",
   "0111001010111101000010111001110011101001001100011111",
   "0111001011110110011110000111110010111101010101101111",
   "0111001100110000000000100001101000110000001101000110",
   "0111001101101001101010001000001110100100001100011111",
   "0111001110100011011010111100011110000010111010100101",
   "0111001111011101010010111111010000111101001011101100",
   "0111010000010111010010010001100001001011000010101100",
   "0111010001010001011000110100001000101011110001111001",
   "0111010010001011100110101000000001100101111100000001",
   "0111010011000101111011101110000110000111010101000000",
   "0111010100000000011000000111010000100101000011000001",
   "0111010100111010111011110100011011011011011111010010",
   "0111010101110101100110110110100001001110010111000100",
   "0111010110110000011001001110011100101000101100100000",
   "0111010111101011010010111101001000011100110111101001",
   "0111011000100110010100000011011111100100100111001101",
   "0111011001100001011100100010011101000001000001101001",
   "0111011010011100101100011010111011111010100101111111",
   "0111011011011000000011101101110111100001001100110100",
   "0111011100010011100010011100001011001100001001001000",
   "0111011101001111001000100110110010011010001001010011",
   "0111011110001010110110001110101000110001011000000010",
   "0111011111000110101011010100101001111111011101010000",
   "0111100000000010100111111001110001111001011111000100",
   "0111100000111110101011111110111100011100000010101001",
   "0111100001111010110111100101000101101011001101010000",
   "0111100010110111001010101101001001110010100101000111",
   "0111100011110011100101011000000101000101010010010111",
   "0111100100110000000111100110110011111110000000000000",
   "0111100101101100110001011010010010111110111100110111",
   "0111100110101001100010110011011110110001111100011111",
   "0111100111100110011011110011010100001000011000001001",
   "0111101000100011011100011010101111111011001111110000",
   "0111101001100000100100101010101111001011001010110100",
   "0111101010011101110100100100001111000000011001011011",
   "0111101011011011001100001000001100101010110101001000",
   "0111101100011000101011010111100101100010000001111111",
   "0111101101010110010010010011010111000101001111011101",
   "0111101110010100000000111100011110111011011001011010",
   "0111101111010001110111010011111010110011001001000010",
   "0111110000001111110101011010101000100010110101110110",
   "0111110001001101111011010001100110001000100110101001",
   "0111110010001100001000111001110001101010010010011111",
   "0111110011001010011110010100001001010101100001100111",
   "0111110100001000111011100001101011011111101110011110",
   "0111110101000111100000100011010110100110000110101101",
   "0111110110000110001101011010001001001101101100000010",
   "0111110111000101000010000111000010000011010101010111",
   "0111111000000011111110101010111111111011101111101001",
   "0111111001000011000011000111000001110011011110111011",
   "0111111010000010001111011100000110101110111111010101",
   "0111111011000001100011101011001101111010100110000000",
   "0111111100000000111111110101010110101010100010001001",
   "0111111101000000100011111011100000011010111101111111",
   "0111111110000000001111111110101010101111111111101111",
   "0111111111000000000011111111110101010101101010101010",
      others => (others => '0'));
      	begin 
      return tmp;
      end init_rom;
	signal rom : memory_t := init_rom;
   signal Y0 :  std_logic_vector(51 downto 0);
begin
	process(clk)
   begin
   if(rising_edge(clk)) then
    if(Enable='1') then
   	Y0 <= rom(  TO_INTEGER(unsigned(X))  );
    end if;
   end if;
   end process;
    Y <= Y0;
end architecture;

--------------------------------------------------------------------------------
--                       LeftShifter_48_by_max_58_uid41
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter_48_by_max_58_uid41 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(47 downto 0);
          S : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(105 downto 0)   );
end entity;

architecture arch of LeftShifter_48_by_max_58_uid41 is
signal level0, level0_d1 :  std_logic_vector(47 downto 0);
signal ps, ps_d1, ps_d2 :  std_logic_vector(5 downto 0);
signal level1 :  std_logic_vector(48 downto 0);
signal level2 :  std_logic_vector(50 downto 0);
signal level3 :  std_logic_vector(54 downto 0);
signal level4 :  std_logic_vector(62 downto 0);
signal level5, level5_d1 :  std_logic_vector(78 downto 0);
signal level6 :  std_logic_vector(110 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
          if(Enable='1') then
            level0_d1 <=  level0;
            ps_d1 <=  ps;
            ps_d2 <=  ps_d1;
            level5_d1 <=  level5;
          end if;
         end if;
      end process;
   level0<= X;
   ps<= S;
   ----------------Synchro barrier, entering cycle 1----------------
   level1<= level0_d1 & (0 downto 0 => '0') when ps_d1(0)= '1' else     (0 downto 0 => '0') & level0_d1;
   level2<= level1 & (1 downto 0 => '0') when ps_d1(1)= '1' else     (1 downto 0 => '0') & level1;
   level3<= level2 & (3 downto 0 => '0') when ps_d1(2)= '1' else     (3 downto 0 => '0') & level2;
   level4<= level3 & (7 downto 0 => '0') when ps_d1(3)= '1' else     (7 downto 0 => '0') & level3;
   level5<= level4 & (15 downto 0 => '0') when ps_d1(4)= '1' else     (15 downto 0 => '0') & level4;
   ----------------Synchro barrier, entering cycle 2----------------
   level6<= level5_d1 & (31 downto 0 => '0') when ps_d2(5)= '1' else     (31 downto 0 => '0') & level5_d1;
   R <= level6(105 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_75_f400_uid127
--                     (IntAdderClassical_75_f400_uid129)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_75_f400_uid127 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(74 downto 0);
          Y : in  std_logic_vector(74 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(74 downto 0)   );
end entity;

architecture arch of IntAdder_75_f400_uid127 is
signal x0 :  std_logic_vector(41 downto 0);
signal y0 :  std_logic_vector(41 downto 0);
signal x1, x1_d1 :  std_logic_vector(32 downto 0);
signal y1, y1_d1 :  std_logic_vector(32 downto 0);
signal sum0, sum0_d1 :  std_logic_vector(42 downto 0);
signal sum1 :  std_logic_vector(33 downto 0);
signal X_d1 :  std_logic_vector(74 downto 0);
signal Y_d1 :  std_logic_vector(74 downto 0);
signal Cin_d1 : std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
          if(Enable='1') then
            x1_d1 <=  x1;
            y1_d1 <=  y1;
            sum0_d1 <=  sum0;
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
          end if;
         end if;
      end process;
   --Classical
   ----------------Synchro barrier, entering cycle 1----------------
   x0 <= X_d1(41 downto 0);
   y0 <= Y_d1(41 downto 0);
   x1 <= X_d1(74 downto 42);
   y1 <= Y_d1(74 downto 42);
   sum0 <= ( "0" & x0) + ( "0" & y0)  + Cin_d1;
   ----------------Synchro barrier, entering cycle 2----------------
   sum1 <= ( "0" & x1_d1) + ( "0" & y1_d1)  + sum0_d1(42);
   R <= sum1(32 downto 0) & sum0_d1(41 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiAdder_75_op2_f400_uid123
--                      (IntCompressorTree_75_2_uid125)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2009-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiAdder_75_op2_f400_uid123 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X0 : in  std_logic_vector(74 downto 0);
          X1 : in  std_logic_vector(74 downto 0);
          R : out  std_logic_vector(74 downto 0)   );
end entity;

architecture arch of IntMultiAdder_75_op2_f400_uid123 is
   component IntAdder_75_f400_uid127 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL , rst : in std_logic;
             X : in  std_logic_vector(74 downto 0);
             Y : in  std_logic_vector(74 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(74 downto 0)   );
   end component;

signal l_0_s_0 :  std_logic_vector(74 downto 0);
signal l_0_s_1 :  std_logic_vector(74 downto 0);
signal myR :  std_logic_vector(74 downto 0);
begin
   l_0_s_0 <= X0;
   l_0_s_1 <= X1;
   FinalAdder_CompressorTree: IntAdder_75_f400_uid127  -- pipelineDepth=2 maxInDelay=2.40572e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 Cin => '0',
                 R => myR,
                 X => l_0_s_0,
                 Y => l_0_s_1);

   ----------------Synchro barrier, entering cycle 2----------------
   R <= myR;
 -- delay at adder output 1.427e-09
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplier_42_43_unsigned_uid119
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Sebastian Banescu (2008-2009)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library work;
entity IntMultiplier_42_43_unsigned_uid119 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(41 downto 0);
          Y : in  std_logic_vector(42 downto 0);
          R : out  std_logic_vector(84 downto 0)   );
end entity;

architecture arch of IntMultiplier_42_43_unsigned_uid119 is
   component IntMultiAdder_75_op2_f400_uid123 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             X0 : in  std_logic_vector(74 downto 0);
             X1 : in  std_logic_vector(74 downto 0);
             R : out  std_logic_vector(74 downto 0)   );
   end component;

signal sX :  std_logic_vector(47 downto 0);
signal sY :  std_logic_vector(50 downto 0);
signal x0, x0_d1, x0_d2, x0_d3 :  std_logic_vector(23 downto 0);
signal x1, x1_d1, x1_d2, x1_d3 :  std_logic_vector(23 downto 0);
signal y0, y0_d1 :  std_logic_vector(16 downto 0);
signal y1, y1_d1, y1_d2 :  std_logic_vector(16 downto 0);
signal y2, y2_d1, y2_d2, y2_d3 :  std_logic_vector(16 downto 0);
signal px0y0, px0y0_d1, px0y0_d2, px0y0_d3 :  std_logic_vector(40 downto 0);
signal tpx0y1 :  std_logic_vector(40 downto 0);
signal px0y1, px0y1_d1, px0y1_d2 :  std_logic_vector(41 downto 0);
signal tpx0y2 :  std_logic_vector(40 downto 0);
signal px0y2, px0y2_d1 :  std_logic_vector(41 downto 0);
signal px1y0, px1y0_d1, px1y0_d2, px1y0_d3 :  std_logic_vector(40 downto 0);
signal tpx1y1 :  std_logic_vector(40 downto 0);
signal px1y1, px1y1_d1, px1y1_d2 :  std_logic_vector(41 downto 0);
signal tpx1y2 :  std_logic_vector(40 downto 0);
signal px1y2, px1y2_d1 :  std_logic_vector(41 downto 0);
signal sum0 :  std_logic_vector(74 downto 0);
signal sum1 :  std_logic_vector(74 downto 0);
signal sum0Low, sum0Low_d1, sum0Low_d2 :  std_logic_vector(23 downto 0);
signal addOp0 :  std_logic_vector(74 downto 0);
signal addOp1 :  std_logic_vector(74 downto 0);
signal addRes :  std_logic_vector(74 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
          if(Enable='1') then
            x0_d1 <=  x0;
            x0_d2 <=  x0_d1;
            x0_d3 <=  x0_d2;
            x1_d1 <=  x1;
            x1_d2 <=  x1_d1;
            x1_d3 <=  x1_d2;
            y0_d1 <=  y0;
            y1_d1 <=  y1;
            y1_d2 <=  y1_d1;
            y2_d1 <=  y2;
            y2_d2 <=  y2_d1;
            y2_d3 <=  y2_d2;
            px0y0_d1 <=  px0y0;
            px0y0_d2 <=  px0y0_d1;
            px0y0_d3 <=  px0y0_d2;
            px0y1_d1 <=  px0y1;
            px0y1_d2 <=  px0y1_d1;
            px0y2_d1 <=  px0y2;
            px1y0_d1 <=  px1y0;
            px1y0_d2 <=  px1y0_d1;
            px1y0_d3 <=  px1y0_d2;
            px1y1_d1 <=  px1y1;
            px1y1_d2 <=  px1y1_d1;
            px1y2_d1 <=  px1y2;
            sum0Low_d1 <=  sum0Low;
            sum0Low_d2 <=  sum0Low_d1;
          end if;
         end if;
      end process;
   sX <= X & "000000";
   sY <= Y & "00000000";
   x0 <= sX(23 downto 0);
   x1 <= sX(47 downto 24);
   y0 <= sY(16 downto 0);
   y1 <= sY(33 downto 17);
   y2 <= sY(50 downto 34);
   ----------------Synchro barrier, entering cycle 1----------------
   px0y0 <= x0_d1 * y0_d1;
   ----------------Synchro barrier, entering cycle 2----------------
   tpx0y1 <= x0_d2 * y1_d2;
   px0y1 <= ( "0" & tpx0y1) + px0y0_d1(40 downto 17);
   ----------------Synchro barrier, entering cycle 3----------------
   tpx0y2 <= x0_d3 * y2_d3;
   px0y2 <= ( "0" & tpx0y2) + px0y1_d1(40 downto 17);
   ----------------Synchro barrier, entering cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   px1y0 <= x1_d1 * y0_d1;
   ----------------Synchro barrier, entering cycle 2----------------
   tpx1y1 <= x1_d2 * y1_d2;
   px1y1 <= ( "0" & tpx1y1) + px1y0_d1(40 downto 17);
   ----------------Synchro barrier, entering cycle 3----------------
   tpx1y2 <= x1_d3 * y2_d3;
   px1y2 <= ( "0" & tpx1y2) + px1y1_d1(40 downto 17);
   ----------------Synchro barrier, entering cycle 4----------------
   sum0 <= px0y2_d1(40 downto 0) & px0y1_d2(16 downto 0) & px0y0_d3(16 downto 0);
   sum1 <= px1y2_d1(40 downto 0) & px1y1_d2(16 downto 0) & px1y0_d3(16 downto 0);
   sum0Low <= sum0(23 downto 0);
   addOp0 <= "000000000000000000000000" & sum0(74 downto 24);
   addOp1 <= "" & sum1(74 downto 0);
   adder: IntMultiAdder_75_op2_f400_uid123  -- pipelineDepth=2 maxInDelay=1.961e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                  rst  => rst,
                 R => addRes,
                 X0 => addOp0,
                 X1 => addOp1);
   ----------------Synchro barrier, entering cycle 6----------------
   R <= addRes(74 downto 0) & sum0Low_d2(23 downto 14);
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_57_f400_uid139
--                     (IntAdderClassical_57_f400_uid141)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_57_f400_uid139 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(56 downto 0);
          Y : in  std_logic_vector(56 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(56 downto 0)   );
end entity;

architecture arch of IntAdder_57_f400_uid139 is
signal x0 :  std_logic_vector(41 downto 0);
signal y0 :  std_logic_vector(41 downto 0);
signal x1, x1_d1 :  std_logic_vector(14 downto 0);
signal y1, y1_d1 :  std_logic_vector(14 downto 0);
signal sum0, sum0_d1 :  std_logic_vector(42 downto 0);
signal sum1 :  std_logic_vector(15 downto 0);
signal X_d1 :  std_logic_vector(56 downto 0);
signal Y_d1 :  std_logic_vector(56 downto 0);
signal Cin_d1 : std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
          if(Enable='1') then
            x1_d1 <=  x1;
            y1_d1 <=  y1;
            sum0_d1 <=  sum0;
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
          end if;
         end if;
      end process;
   --Classical
   ----------------Synchro barrier, entering cycle 1----------------
   x0 <= X_d1(41 downto 0);
   y0 <= Y_d1(41 downto 0);
   x1 <= X_d1(56 downto 42);
   y1 <= Y_d1(56 downto 42);
   sum0 <= ( "0" & x0) + ( "0" & y0)  + Cin_d1;
   ----------------Synchro barrier, entering cycle 2----------------
   sum1 <= ( "0" & x1_d1) + ( "0" & y1_d1)  + sum0_d1(42);
   R <= sum1(14 downto 0) & sum0_d1(41 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_52_f400_uid133
--                     (IntAdderClassical_52_f400_uid135)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_52_f400_uid133 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(51 downto 0);
          Y : in  std_logic_vector(51 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(51 downto 0)   );
end entity;

architecture arch of IntAdder_52_f400_uid133 is
signal x0 :  std_logic_vector(41 downto 0);
signal y0 :  std_logic_vector(41 downto 0);
signal x1, x1_d1 :  std_logic_vector(9 downto 0);
signal y1, y1_d1 :  std_logic_vector(9 downto 0);
signal sum0, sum0_d1 :  std_logic_vector(42 downto 0);
signal sum1 :  std_logic_vector(10 downto 0);
signal X_d1 :  std_logic_vector(51 downto 0);
signal Y_d1 :  std_logic_vector(51 downto 0);
signal Cin_d1 : std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
          if(Enable='1') then
            x1_d1 <=  x1;
            y1_d1 <=  y1;
            sum0_d1 <=  sum0;
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
          end if;
         end if;
      end process;
   --Classical
   ----------------Synchro barrier, entering cycle 1----------------
   x0 <= X_d1(41 downto 0);
   y0 <= Y_d1(41 downto 0);
   x1 <= X_d1(51 downto 42);
   y1 <= Y_d1(51 downto 42);
   sum0 <= ( "0" & x0) + ( "0" & y0)  + Cin_d1;
   ----------------Synchro barrier, entering cycle 2----------------
   sum1 <= ( "0" & x1_d1) + ( "0" & y1_d1)  + sum0_d1(42);
   R <= sum1(9 downto 0) & sum0_d1(41 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_51_f484_uid61
--                     (IntAdderClassical_51_f484_uid63)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_51_f484_uid61 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(50 downto 0);
          Y : in  std_logic_vector(50 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(50 downto 0)   );
end entity;

architecture arch of IntAdder_51_f484_uid61 is
signal x0 :  std_logic_vector(22 downto 0);
signal y0 :  std_logic_vector(22 downto 0);
signal x1, x1_d1 :  std_logic_vector(22 downto 0);
signal y1, y1_d1 :  std_logic_vector(22 downto 0);
signal x2, x2_d1, x2_d2 :  std_logic_vector(4 downto 0);
signal y2, y2_d1, y2_d2 :  std_logic_vector(4 downto 0);
signal sum0, sum0_d1, sum0_d2 :  std_logic_vector(23 downto 0);
signal sum1, sum1_d1 :  std_logic_vector(23 downto 0);
signal sum2 :  std_logic_vector(5 downto 0);
signal X_d1 :  std_logic_vector(50 downto 0);
signal Y_d1 :  std_logic_vector(50 downto 0);
signal Cin_d1 : std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
          if(Enable='1') then
            x1_d1 <=  x1;
            y1_d1 <=  y1;
            x2_d1 <=  x2;
            x2_d2 <=  x2_d1;
            y2_d1 <=  y2;
            y2_d2 <=  y2_d1;
            sum0_d1 <=  sum0;
            sum0_d2 <=  sum0_d1;
            sum1_d1 <=  sum1;
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
          end if;
         end if;
      end process;
   --Classical
   ----------------Synchro barrier, entering cycle 1----------------
   x0 <= X_d1(22 downto 0);
   y0 <= Y_d1(22 downto 0);
   x1 <= X_d1(45 downto 23);
   y1 <= Y_d1(45 downto 23);
   x2 <= X_d1(50 downto 46);
   y2 <= Y_d1(50 downto 46);
   sum0 <= ( "0" & x0) + ( "0" & y0)  + Cin_d1;
   ----------------Synchro barrier, entering cycle 2----------------
   sum1 <= ( "0" & x1_d1) + ( "0" & y1_d1)  + sum0_d1(23);
   ----------------Synchro barrier, entering cycle 3----------------
   sum2 <= ( "0" & x2_d2) + ( "0" & y2_d2)  + sum1_d1(23);
   R <= sum2(4 downto 0) & sum1_d1(22 downto 0) & sum0_d2(22 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_43_f400_uid113
--                     (IntAdderClassical_43_f400_uid115)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_43_f400_uid113 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL , rst : in std_logic;
          X : in  std_logic_vector(42 downto 0);
          Y : in  std_logic_vector(42 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(42 downto 0)   );
end entity;

architecture arch of IntAdder_43_f400_uid113 is
signal x0 :  std_logic_vector(41 downto 0);
signal y0 :  std_logic_vector(41 downto 0);
signal x1, x1_d1 :  std_logic_vector(0 downto 0);
signal y1, y1_d1 :  std_logic_vector(0 downto 0);
signal sum0, sum0_d1 :  std_logic_vector(42 downto 0);
signal sum1 :  std_logic_vector(1 downto 0);
signal X_d1 :  std_logic_vector(42 downto 0);
signal Y_d1 :  std_logic_vector(42 downto 0);
signal Cin_d1 : std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
          if(Enable='1') then
            x1_d1 <=  x1;
            y1_d1 <=  y1;
            sum0_d1 <=  sum0;
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
           end if;
         end if;
      end process;
   --Classical
   ----------------Synchro barrier, entering cycle 1----------------
   x0 <= X_d1(41 downto 0);
   y0 <= Y_d1(41 downto 0);
   x1 <= X_d1(42 downto 42);
   y1 <= Y_d1(42 downto 42);
   sum0 <= ( "0" & x0) + ( "0" & y0)  + Cin_d1;
   ----------------Synchro barrier, entering cycle 2----------------
   sum1 <= ( "0" & x1_d1) + ( "0" & y1_d1)  + sum0_d1(42);
   R <= sum1(0 downto 0) & sum0_d1(41 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_43_f400_uid107
--                     (IntAdderClassical_43_f400_uid109)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_43_f400_uid107 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(42 downto 0);
          Y : in  std_logic_vector(42 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(42 downto 0)   );
end entity;

architecture arch of IntAdder_43_f400_uid107 is
signal x0 :  std_logic_vector(41 downto 0);
signal y0 :  std_logic_vector(41 downto 0);
signal x1, x1_d1 :  std_logic_vector(0 downto 0);
signal y1, y1_d1 :  std_logic_vector(0 downto 0);
signal sum0, sum0_d1 :  std_logic_vector(42 downto 0);
signal sum1 :  std_logic_vector(1 downto 0);
signal X_d1 :  std_logic_vector(42 downto 0);
signal Y_d1 :  std_logic_vector(42 downto 0);
signal Cin_d1 : std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
          if(Enable='1') then
            x1_d1 <=  x1;
            y1_d1 <=  y1;
            sum0_d1 <=  sum0;
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
          end if;
         end if;
      end process;
   --Classical
   ----------------Synchro barrier, entering cycle 1----------------
   x0 <= X_d1(41 downto 0);
   y0 <= Y_d1(41 downto 0);
   x1 <= X_d1(42 downto 42);
   y1 <= Y_d1(42 downto 42);
   sum0 <= ( "0" & x0) + ( "0" & y0)  + Cin_d1;
   ----------------Synchro barrier, entering cycle 2----------------
   sum1 <= ( "0" & x1_d1) + ( "0" & y1_d1)  + sum0_d1(42);
   R <= sum1(0 downto 0) & sum0_d1(41 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_56_f400_uid95
--                    (IntAdderAlternative_56_f400_uid99)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_56_f400_uid95 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(55 downto 0);
          Y : in  std_logic_vector(55 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(55 downto 0)   );
end entity;

architecture arch of IntAdder_56_f400_uid95 is
signal s_sum_l0_idx0 :  std_logic_vector(40 downto 0);
signal s_sum_l0_idx1, s_sum_l0_idx1_d1 :  std_logic_vector(16 downto 0);
signal sum_l0_idx0, sum_l0_idx0_d1 :  std_logic_vector(39 downto 0);
signal c_l0_idx0, c_l0_idx0_d1 :  std_logic_vector(0 downto 0);
signal sum_l0_idx1 :  std_logic_vector(15 downto 0);
signal c_l0_idx1 :  std_logic_vector(0 downto 0);
signal s_sum_l1_idx1 :  std_logic_vector(16 downto 0);
signal sum_l1_idx1 :  std_logic_vector(15 downto 0);
signal c_l1_idx1 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
           if(Enable='1') then
            s_sum_l0_idx1_d1 <=  s_sum_l0_idx1;
            sum_l0_idx0_d1 <=  sum_l0_idx0;
            c_l0_idx0_d1 <=  c_l0_idx0;
           end if;
         end if;
      end process;
   --Alternative
   s_sum_l0_idx0 <= ( "0" & X(39 downto 0)) + ( "0" & Y(39 downto 0)) + Cin;
   s_sum_l0_idx1 <= ( "0" & X(55 downto 40)) + ( "0" & Y(55 downto 40));
   sum_l0_idx0 <= s_sum_l0_idx0(39 downto 0);
   c_l0_idx0 <= s_sum_l0_idx0(40 downto 40);
   sum_l0_idx1 <= s_sum_l0_idx1(15 downto 0);
   c_l0_idx1 <= s_sum_l0_idx1(16 downto 16);
   ----------------Synchro barrier, entering cycle 1----------------
   s_sum_l1_idx1 <=  s_sum_l0_idx1_d1 + c_l0_idx0_d1(0 downto 0);
   sum_l1_idx1 <= s_sum_l1_idx1(15 downto 0);
   c_l1_idx1 <= s_sum_l1_idx1(16 downto 16);
   R <= sum_l1_idx1(15 downto 0) & sum_l0_idx0_d1(39 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiAdder_56_op2_f400_uid91
--                       (IntCompressorTree_56_2_uid93)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2009-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiAdder_56_op2_f400_uid91 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X0 : in  std_logic_vector(55 downto 0);
          X1 : in  std_logic_vector(55 downto 0);
          R : out  std_logic_vector(55 downto 0)   );
end entity;

architecture arch of IntMultiAdder_56_op2_f400_uid91 is
   component IntAdder_56_f400_uid95 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             X : in  std_logic_vector(55 downto 0);
             Y : in  std_logic_vector(55 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(55 downto 0)   );
   end component;

signal l_0_s_0 :  std_logic_vector(55 downto 0);
signal l_0_s_1 :  std_logic_vector(55 downto 0);
signal myR :  std_logic_vector(55 downto 0);
begin
   l_0_s_0 <= X0;
   l_0_s_1 <= X1;
   FinalAdder_CompressorTree: IntAdder_56_f400_uid95  -- pipelineDepth=1 maxInDelay=8.8944e-10
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 Cin => '0',
                 R => myR,
                 X => l_0_s_0,
                 Y => l_0_s_1);

   ----------------Synchro barrier, entering cycle 1----------------
   R <= myR;
 -- delay at adder output 1.036e-09
end architecture;

--------------------------------------------------------------------------------
--                     IntTruncMultiplier_26_31_31_signed
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Sebastian Banescu, Bogdan Pasca, Radu Tudoran (2010-2011)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
library work;
entity IntTruncMultiplier_26_31_31_signed is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(25 downto 0);
          Y : in  std_logic_vector(30 downto 0);
          R_old : out  std_logic_vector(30 downto 0);
          R : out  std_logic_vector(30 downto 0)   );
end entity;

architecture arch of IntTruncMultiplier_26_31_31_signed is
   component IntMultiAdder_56_op2_f400_uid91 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             X0 : in  std_logic_vector(55 downto 0);
             X1 : in  std_logic_vector(55 downto 0);
             R : out  std_logic_vector(55 downto 0)   );
   end component;

signal x0_0 :  std_logic_vector(24 downto 0);
signal y0_0 :  std_logic_vector(17 downto 0);
signal pxy00 :  std_logic_vector(42 downto 0);
signal addOpDSP0, addOpDSP0_d1, addOpDSP0_d2, addOpDSP0_d3  :  std_logic_vector(55 downto 0);
signal x1_0 :  std_logic_vector(24 downto 0);
signal y1_0 :  std_logic_vector(17 downto 0);
signal pxy10, pxy10_d1, pxy10_d2 :  std_logic_vector(42 downto 0);
signal x1_1, x1_1_d1 :  std_logic_vector(24 downto 0);
signal y1_1, y1_1_d1 :  std_logic_vector(17 downto 0);
signal txy11 :  std_logic_vector(42 downto 0);
signal pxy11, pxy11_d1 :  std_logic_vector(42 downto 0);
signal addOpDSP1, addOpDSP1_d1 :  std_logic_vector(55 downto 0);
signal addRes :  std_logic_vector(55 downto 0);

signal addResOld :  std_logic_vector(55 downto 0);

begin
   process(clk)
      begin
         if clk'event and clk = '1' then
           if(Enable='1') then
            addOpDSP0_d1 <=  addOpDSP0;
            addOpDSP0_d2 <=  addOpDSP0_d1;
            addOpDSP0_d3 <=  addOpDSP0_d2;
            addOpDSP1_d1 <=  addOpDSP1   ;
            pxy10_d1 <=  pxy10;
            pxy10_d2 <=  pxy10_d1;
            x1_1_d1 <=  x1_1;
            y1_1_d1 <=  y1_1;
            pxy11_d1 <=  pxy11;
           end if;
         end if;
      end process;
   ----------------Synchro barrier, entering cycle 0----------------
   ----------------Synchro barrier, entering cycle 0----------------
   x0_0 <= "0" & "" & X(0 downto 0) & "00000000000000000000000";
   y0_0 <="" & Y(30 downto 13) & "";
   pxy00 <= x0_0(24 downto 0) * y0_0(17 downto 0); --0
   addOpDSP0 <= (25 downto 0 => pxy00(40)) & pxy00(40 downto 23) & "000000000000"; --1
   ----------------Synchro barrier, entering cycle 0----------------
   ----------------Synchro barrier, entering cycle 0----------------
   x1_0 <= "" & X(25 downto 1) & "";
   y1_0 <= "0" & "" & Y(12 downto 0) & "0000";
   pxy10 <= x1_0(24 downto 0) * y1_0(17 downto 0); --0
   ----------------Synchro barrier, entering cycle 0----------------
   x1_1 <= "" & X(25 downto 1) & "";
   y1_1 <="" & Y(30 downto 13) & "";
   ----------------Synchro barrier, entering cycle 1----------------
   txy11 <= x1_1_d1(24 downto 0) * y1_1_d1(17 downto 0);
   pxy11 <= (txy11(42 downto 0)) + ((16 downto 0 => pxy10_d1(42)) &pxy10_d1(42 downto 17));
   ----------------Synchro barrier, entering cycle 2----------------
   addOpDSP1 <= (0 downto 0 => pxy11_d1(41)) & pxy11_d1(41 downto 0) & pxy10_d2(16 downto 4) & "" &  "";--3 bpadX 0 bpadY 4
   adder: IntMultiAdder_56_op2_f400_uid91  -- pipelineDepth=1 maxInDelay=4.4472e-10
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 R => addRes,
                 X0 => addOpDSP0_d3,  -- +1 CHGMNT OF
                 X1 => addOpDSP1_d1); -- +1 CHGMNT OF

   adder2: IntMultiAdder_56_op2_f400_uid91  -- pipelineDepth=1 maxInDelay=4.4472e-10
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 R => addResOld,
                 X0 => addOpDSP0_d2, 
                 X1 => addOpDSP1); 

   ----------------Synchro barrier, entering cycle 3----------------
   R_old <= addResOld(55 downto 25);
   R <= addRes(55 downto 25);
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_48_f400_uid78
--                    (IntAdderAlternative_48_f400_uid82)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_48_f400_uid78 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(47 downto 0);
          Y : in  std_logic_vector(47 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntAdder_48_f400_uid78 is
signal s_sum_l0_idx0 :  std_logic_vector(40 downto 0);
signal s_sum_l0_idx1, s_sum_l0_idx1_d1 :  std_logic_vector(8 downto 0);
signal sum_l0_idx0, sum_l0_idx0_d1 :  std_logic_vector(39 downto 0);
signal c_l0_idx0, c_l0_idx0_d1 :  std_logic_vector(0 downto 0);
signal sum_l0_idx1 :  std_logic_vector(7 downto 0);
signal c_l0_idx1 :  std_logic_vector(0 downto 0);
signal s_sum_l1_idx1 :  std_logic_vector(8 downto 0);
signal sum_l1_idx1 :  std_logic_vector(7 downto 0);
signal c_l1_idx1 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
           if(Enable='1') then
            s_sum_l0_idx1_d1 <=  s_sum_l0_idx1;
            sum_l0_idx0_d1 <=  sum_l0_idx0;
            c_l0_idx0_d1 <=  c_l0_idx0;
           end if;
         end if;
      end process;
   --Alternative
   s_sum_l0_idx0 <= ( "0" & X(39 downto 0)) + ( "0" & Y(39 downto 0)) + Cin;
   s_sum_l0_idx1 <= ( "0" & X(47 downto 40)) + ( "0" & Y(47 downto 40));
   sum_l0_idx0 <= s_sum_l0_idx0(39 downto 0);
   c_l0_idx0 <= s_sum_l0_idx0(40 downto 40);
   sum_l0_idx1 <= s_sum_l0_idx1(7 downto 0);
   c_l0_idx1 <= s_sum_l0_idx1(8 downto 8);
   ----------------Synchro barrier, entering cycle 1----------------
   s_sum_l1_idx1 <=  s_sum_l0_idx1_d1 + c_l0_idx0_d1(0 downto 0);
   sum_l1_idx1 <= s_sum_l1_idx1(7 downto 0);
   c_l1_idx1 <= s_sum_l1_idx1(8 downto 8);
   R <= sum_l1_idx1(7 downto 0) & sum_l0_idx0_d1(39 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                      IntMultiAdder_48_op2_f400_uid74
--                       (IntCompressorTree_48_2_uid76)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2009-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiAdder_48_op2_f400_uid74 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X0 : in  std_logic_vector(47 downto 0);
          X1 : in  std_logic_vector(47 downto 0);
          R : out  std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiAdder_48_op2_f400_uid74 is
   component IntAdder_48_f400_uid78 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             X : in  std_logic_vector(47 downto 0);
             Y : in  std_logic_vector(47 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(47 downto 0)   );
   end component;

signal l_0_s_0 :  std_logic_vector(47 downto 0);
signal l_0_s_1 :  std_logic_vector(47 downto 0);
signal myR :  std_logic_vector(47 downto 0);
begin
   l_0_s_0 <= X0;
   l_0_s_1 <= X1;
   FinalAdder_CompressorTree: IntAdder_48_f400_uid78  -- pipelineDepth=1 maxInDelay=8.8944e-10
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 Cin => '0',
                 R => myR,
                 X => l_0_s_0,
                 Y => l_0_s_1);

   ----------------Synchro barrier, entering cycle 1----------------
   R <= myR;
 -- delay at adder output 8.52e-10
end architecture;
--------------------------------------------------------------------------------
--                     IntTruncMultiplier_25_23_23_signed
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Sebastian Banescu, Bogdan Pasca, Radu Tudoran (2010-2011)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
library work;
entity IntTruncMultiplier_25_23_23_signed is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(24 downto 0);
          Y : in  std_logic_vector(22 downto 0);
          R : out  std_logic_vector(22 downto 0)   );
end entity;

architecture arch of IntTruncMultiplier_25_23_23_signed is
   component IntMultiAdder_48_op2_f400_uid74 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OF, rst : in std_logic;
             X0 : in  std_logic_vector(47 downto 0);
             X1 : in  std_logic_vector(47 downto 0);
             R : out  std_logic_vector(47 downto 0)   );
   end component;

signal x0_0 :  std_logic_vector(24 downto 0);
signal y0_0 :  std_logic_vector(17 downto 0);
signal pxy00, pxy00_d1, pxy00_d2 :  std_logic_vector(42 downto 0);
signal x0_1, x0_1_d1 :  std_logic_vector(24 downto 0);
signal y0_1, y0_1_d1 :  std_logic_vector(17 downto 0);
signal txy01 :  std_logic_vector(42 downto 0);
signal pxy01, pxy01_d1 :  std_logic_vector(42 downto 0);
signal addOpDSP0 :  std_logic_vector(47 downto 0);
signal addRes :  std_logic_vector(47 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
           if(Enable='1') then
            pxy00_d1 <=  pxy00;
            pxy00_d2 <=  pxy00_d1;
            x0_1_d1 <=  x0_1;
            y0_1_d1 <=  y0_1;
            pxy01_d1 <=  pxy01;
           end if;
         end if;
      end process;
   ----------------Synchro barrier, entering cycle 0----------------
   ----------------Synchro barrier, entering cycle 0----------------
   x0_0 <= "" & X(24 downto 0) & "";
   y0_0 <= "0" & "" & Y(4 downto 0) & "000000000000";
   pxy00 <= x0_0(24 downto 0) * y0_0(17 downto 0); --0
   ----------------Synchro barrier, entering cycle 0----------------
   x0_1 <= "" & X(24 downto 0) & "";
   y0_1 <="" & Y(22 downto 5) & "";
   ----------------Synchro barrier, entering cycle 1----------------
   txy01 <= x0_1_d1(24 downto 0) * y0_1_d1(17 downto 0);
   pxy01 <= (txy01(42 downto 0)) + ((16 downto 0 => pxy00_d1(42)) &pxy00_d1(42 downto 17));
   ----------------Synchro barrier, entering cycle 2----------------
   addOpDSP0 <= (0 downto 0 => pxy01_d1(41)) & pxy01_d1(41 downto 0) & pxy00_d2(16 downto 12) & "" &  "";--3 bpadX 0 bpadY 12
   adder: IntMultiAdder_48_op2_f400_uid74  -- pipelineDepth=1 maxInDelay=4.4472e-10
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 R => addRes,
                 X0 => addOpDSP0,
                 X1 => "000000000000000000000010000000000000000000000000");
   ----------------Synchro barrier, entering cycle 3----------------
   R <= addRes(47 downto 25);
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_37_f400_uid101
--                     (IntAdderClassical_37_f400_uid103)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_37_f400_uid101 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL , rst : in std_logic;
          X : in  std_logic_vector(36 downto 0);
          Y : in  std_logic_vector(36 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(36 downto 0)   );
end entity;

architecture arch of IntAdder_37_f400_uid101 is
signal X_d1 :  std_logic_vector(36 downto 0);
signal Y_d1 :  std_logic_vector(36 downto 0);
signal Cin_d1 : std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
           if(Enable='1') then
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
           end if;
         end if;
      end process;
   --Classical
   ----------------Synchro barrier, entering cycle 1----------------
    R <= X_d1 + Y_d1 + Cin_d1;
end architecture;
--------------------------------------------------------------------------------
--                           IntAdder_31_f400_uid84
--                    (IntAdderAlternative_31_f400_uid88)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_31_f400_uid84 is
   port (-- OL clk, rst : in std_logic;
          X : in  std_logic_vector(30 downto 0);
          Y : in  std_logic_vector(30 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(30 downto 0)   );
end entity;

architecture arch of IntAdder_31_f400_uid84 is
begin
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                     PolynomialEvaluator_degree2_uid71
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity PolynomialEvaluator_degree2_uid71 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          Y : in  std_logic_vector(24 downto 0);
          a0 : in  std_logic_vector(35 downto 0);
          a1 : in  std_logic_vector(29 downto 0);
          a2 : in  std_logic_vector(22 downto 0);
          R_old : out  std_logic_vector(36 downto 0);
          R : out  std_logic_vector(36 downto 0)   );
end entity;

architecture arch of PolynomialEvaluator_degree2_uid71 is
   component IntAdder_31_f400_uid84 is
      port ( -- OL clk : in std_logic;
             -- OL Enable : in std_logic;
-- OL,, rst : in std_logic;
             X : in  std_logic_vector(30 downto 0);
             Y : in  std_logic_vector(30 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(30 downto 0)   );
   end component;

   component IntAdder_37_f400_uid101 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL,, rst : in std_logic;
             X : in  std_logic_vector(36 downto 0);
             Y : in  std_logic_vector(36 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(36 downto 0)   );
   end component;

   component IntTruncMultiplier_25_23_23_signed is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL,, rst : in std_logic;
             X : in  std_logic_vector(24 downto 0);
             Y : in  std_logic_vector(22 downto 0);
             R : out  std_logic_vector(22 downto 0)   );
   end component;

   component IntTruncMultiplier_26_31_31_signed is
      port ( clk  : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             X : in  std_logic_vector(25 downto 0);
             Y : in  std_logic_vector(30 downto 0);
             R_old : out  std_logic_vector(30 downto 0);
             R : out  std_logic_vector(30 downto 0)   );
   end component;

signal sigmaP0, sigmaP0_d1 :  std_logic_vector(22 downto 0);
signal yT1, yT1_d1 :  std_logic_vector(24 downto 0);
signal piPT1 :  std_logic_vector(22 downto 0);
signal op1_1 :  std_logic_vector(30 downto 0);
signal op2_1 :  std_logic_vector(30 downto 0);
signal sigmaP1 :  std_logic_vector(30 downto 0);
signal yT2 :  std_logic_vector(25 downto 0);
signal piP2 :  std_logic_vector(30 downto 0);
signal piP2_old :  std_logic_vector(30 downto 0);
signal op1_2_old :  std_logic_vector(36 downto 0);
signal op2_2_old :  std_logic_vector(36 downto 0);
signal op1_2 :  std_logic_vector(36 downto 0);
signal op2_2 :  std_logic_vector(36 downto 0);
signal sigmaP2_old :  std_logic_vector(36 downto 0);
signal sigmaP2 :  std_logic_vector(36 downto 0);
signal Y_d1, Y_d2, Y_d3, Y_d4 :  std_logic_vector(24 downto 0);
signal a0_d1, a0_d2, a0_d3, a0_d4, a0_d5, a0_d6, a0_d7, a0_d8 :  std_logic_vector(35 downto 0);
signal a1_d1, a1_d2, a1_d3, a1_d4 :  std_logic_vector(29 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
           if(Enable='1') then
            sigmaP0_d1 <=  sigmaP0;
            yT1_d1 <=  yT1;
            Y_d1 <=  Y;
            Y_d2 <=  Y_d1;
            Y_d3 <=  Y_d2;
            Y_d4 <=  Y_d3;
            a0_d1 <=  a0;
            a0_d2 <=  a0_d1;
            a0_d3 <=  a0_d2;
            a0_d4 <=  a0_d3;
            a0_d5 <=  a0_d4;
            a0_d6 <=  a0_d5;
            a0_d7 <=  a0_d6;
            a0_d8 <=  a0_d7;
            a1_d1 <=  a1;
            a1_d2 <=  a1_d1;
            a1_d3 <=  a1_d2;
            a1_d4 <=  a1_d3;
           end if;
         end if;
      end process;
   -- LSB weight of sigmaP0 is=0 size=23
   sigmaP0 <= a2;
   -- LSB weight of yT1 is=-8 size=25
   yT1 <= "0" & Y(24 downto 1);
   -- LSB weight of piP1 is=-8 size=48
   ----------------Synchro barrier, entering cycle 1----------------
   Product_1: IntTruncMultiplier_25_23_23_signed  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 R => piPT1,
                 X => yT1_d1,
                 Y => sigmaP0_d1);
   ----------------Synchro barrier, entering cycle 4----------------
   op1_1 <= ((0 downto 0 => a1_d4(29)) & a1_d4 & "");
   op2_1 <= ((8 downto 0 => piPT1(21)) & piPT1(21 downto 0) & "");
   Sum1: IntAdder_31_f400_uid84  -- pipelineDepth=0 maxInDelay=8.52e-10
      port map (-- OL clk  => clk,
-- OL                 Enable => Enable,
-- OL                 rst  => rst,
                 Cin => '1',
                 R => sigmaP1,
                 X => op1_1,
                 Y => op2_1);
   -- weight of yT2 is=-8 size=26
   yT2 <= "0" & Y_d4(24 downto 0);
   -- weight of piP2 is=-7 size=57
   Product_2: IntTruncMultiplier_26_31_31_signed  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 R_old => piP2_old,
                 R => piP2,
                 X => yT2,
                 Y => sigmaP1);
   ----------------Synchro barrier, entering cycle 7----------------
   -- the delay at the output of the multiplier is : 1.036e-09
   op1_2_old <= (6 downto 0 => piP2_old(30)) & piP2_old(29 downto 0);
   op1_2 <= (6 downto 0 => piP2(30)) & piP2(29 downto 0);
   op2_2_old <= (0 downto 0 => a0_d7(35)) & a0_d7;
   op2_2 <= (0 downto 0 => a0_d8(35)) & a0_d8; -- + 1 CHGMNT OF
   Sum2: IntAdder_37_f400_uid101  -- pipelineDepth=1 maxInDelay=1.48072e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 Cin => '1',
                 R => sigmaP2,
                 X => op1_2,
                 Y => op2_2);

   Sum22: IntAdder_37_f400_uid101  -- pipelineDepth=1 maxInDelay=1.48072e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 Cin => '1',
                 R => sigmaP2_old,
                 X => op1_2_old,
                 Y => op2_2_old);

   ----------------Synchro barrier, entering cycle 8----------------
   R_old <= sigmaP2_old(36 downto 0);
   R <= sigmaP2(36 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                            PolyCoeffTable_8_89
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Mioara Joldes (2010)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity PolyCoeffTable_8_89 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(7 downto 0);
          Y : out  std_logic_vector(88 downto 0)   );
end entity;

architecture arch of PolyCoeffTable_8_89 is
   -- Build a 2-D array type for the RoM
   subtype word_t is std_logic_vector(44 downto 0);
   type memory_t is array(0 to 511) of word_t;
   function init_rom
      return memory_t is 
      variable tmp : memory_t := (
   "010000000000000000001111111111111111111111111",
   "010000000000000000100100000000010000000000000",
   "010000000000000001011000000000100000000000000",
   "010000000000000001101110000000110000000000000",
   "010000000000000010000100000001000000000000000",
   "010000000000000010111000000001010000000000000",
   "010000000000000011001110000001100000000000001",
   "010000000000000011100100000001110000000000001",
   "010000000000000100011000000010000000000000001",
   "010000000000000100101110000010010000000000010",
   "010000000000000101000100000010100000000000011",
   "010000000000000101110100000010110000000000011",
   "010000000000000110001010000011000000000000100",
   "010000000000000110100110000011010000000000101",
   "010000000000000111010110000011100000000000110",
   "010000000000000111101100000011110000000000111",
   "010000000000001000011100000100000000000000111",
   "010000000000001000110010000100010000000001001",
   "010000000000001001001000000100100000000001010",
   "010000000000001001110100000100110000000001011",
   "010000000000001010010000000101000000000001100",
   "010000000000001010111100000101010000000001101",
   "010000000000001011001110000101100000000001111",
   "010000000000001011100110000101110000000010000",
   "010000000000001100010010000110000000000010001",
   "010000000000001100100110000110010000000010011",
   "010000000000001101010010000110100000000010101",
   "010000000000001101100110000110110000000010110",
   "010000000000001110010100000111000000000011000",
   "010000000000001110111100000111010000000011010",
   "010000000000001111001100000111100000000011100",
   "010000000000001111110110000111110000000011110",
   "010000000000010000001000001000000000000100000",
   "010000000000010000110010001000010000000100010",
   "010000000000010001011000001000100000000100100",
   "010000000000010001111010001000110000000100110",
   "010000000000010010001000001001000000000101000",
   "010000000000010010110000001001010000000101010",
   "010000000000010011001110001001100000000101101",
   "010000000000010011110010001001110000000101111",
   "010000000000010100010010001010000000000110001",
   "010000000000010100110100001010010000000110100",
   "010000000000010101010000001010100000000110111",
   "010000000000010101110010001010110000000111001",
   "010000000000010110001010001011000000000111100",
   "010000000000010110100100001011010000000111111",
   "010000000000010111010100001011100000001000010",
   "010000000000010111110000001011110000001000101",
   "010000000000011000011100001100000000001000111",
   "010000000000011000110000001100010000001001011",
   "010000000000011001011010001100100000001001110",
   "010000000000011001101010001100110000001010001",
   "010000000000011010010010001101000000001010100",
   "010000000000011010111010001101010000001010111",
   "010000000000011011011010001101100000001011011",
   "010000000000011011111010001101110000001011110",
   "010000000000011100010110001110000000001100010",
   "010000000000011100110000001110010000001100101",
   "010000000000011101010000001110100000001101001",
   "010000000000011101111100001110110000001101100",
   "010000000000011110010000001111000000001110000",
   "010000000000011110111010001111010000001110100",
   "010000000000011111001000001111100000001111000",
   "010000000000011111110000001111110000001111100",
   "010000000000100000010000010000000000010000000",
   "010000000000100000101110010000010000010000100",
   "010000000000100001001000010000100000010001000",
   "010000000000100001111000010000110000010001100",
   "010000000000100010001100010001000000010010000",
   "010000000000100010111100010001010000010010100",
   "010000000000100011000110010001100000010011001",
   "010000000000100011101010010001110000010011101",
   "010000000000100100001000010010000000010100010",
   "010000000000100100111100010010010000010100110",
   "010000000000100101010100010010100000010101011",
   "010000000000100101111110010010110000010101111",
   "010000000000100110001100010011000000010110100",
   "010000000000100110101100010011010000010111001",
   "010000000000100111001010010011100000010111110",
   "010000000000100111100110010011110000011000011",
   "010000000000101000010100010100000000011001000",
   "010000000000101001000000010100010000011001101",
   "010000000000101001000110010100100000011010010",
   "010000000000101001101000010100110000011010111",
   "010000000000101010011010010101000000011011100",
   "010000000000101010101110010101010000011100001",
   "010000000000101011010110010101100000011100111",
   "010000000000101011110110010101110000011101100",
   "010000000000101100010010010110000000011110010",
   "010000000000101100101010010110010000011110111",
   "010000000000101101010010010110100000011111101",
   "010000000000101101111000010110110000100000010",
   "010000000000101110010010010111000000100001000",
   "010000000000101110100110010111010000100001110",
   "010000000000101111010010010111100000100010100",
   "010000000000101111110100010111110000100011010",
   "010000000000110000010000011000000000100100000",
   "010000000000110000111010011000010000100100110",
   "010000000000110001001010011000100000100101100",
   "010000000000110001101000011000110000100110010",
   "010000000000110010010110011001000000100111000",
   "010000000000110010101010011001010000100111110",
   "010000000000110011001000011001100000101000101",
   "010000000000110011111010011001110000101001011",
   "010000000000110100001000011010000000101010010",
   "010000000000110100101010011010010000101011000",
   "010000000000110101001000011010100000101011111",
   "010000000000110101110000011010110000101100101",
   "010000000000110110001110011011000000101101100",
   "010000000000110110101000011011010000101110011",
   "010000000000110111001100011011100000101111010",
   "010000000000110111101100011011110000110000001",
   "010000000000111000011100011100000000110001000",
   "010000000000111000101000011100010000110001111",
   "010000000000111001011010011100100000110010110",
   "010000000000111001101110011100110000110011101",
   "010000000000111010001100011101000000110100100",
   "010000000000111010111000011101010000110101011",
   "010000000000111011011110011101100000110110011",
   "010000000000111011111000011101110000110111010",
   "010000000000111100001000011110000000111000010",
   "010000000000111100111110011110010000111001001",
   "010000000000111101001100011110100000111010001",
   "010000000000111101101000011110110000111011000",
   "010000000000111110011010011111000000111100000",
   "010000000000111110111010011111010000111101000",
   "010000000000111111010000011111100000111110000",
   "010000000000111111110000011111110000111111000",
   "010000000001000000100000100000000001000000000",
   "010000000001000000101010100000010001000001000",
   "010000000001000001010110100000100001000010000",
   "010000000001000001110110100000110001000011000",
   "010000000001000010001110100001000001000100000",
   "010000000001000010101110100001010001000101000",
   "010000000001000011010110100001100001000110001",
   "010000000001000011110100100001110001000111001",
   "010000000001000100011110100010000001001000010",
   "010000000001000100111000100010010001001001010",
   "010000000001000101100000100010100001001010011",
   "010000000001000101110010100010110001001011011",
   "010000000001000110011000100011000001001100100",
   "010000000001000110101000100011010001001101101",
   "010000000001000111100000100011100001001110110",
   "010000000001000111101000100011110001001111111",
   "010000000001001000010110100100000001010001000",
   "010000000001001000111000100100010001010010001",
   "010000000001001001001010100100100001010011010",
   "010000000001001001110110100100110001010100011",
   "010000000001001010011000100101000001010101100",
   "010000000001001010100100100101010001010110110",
   "010000000001001011010110100101100001010111111",
   "010000000001001011111000100101110001011001000",
   "010000000001001100100000100110000001011010010",
   "010000000001001100110100100110010001011011011",
   "010000000001001101001110100110100001011100101",
   "010000000001001101110100100110110001011101111",
   "010000000001001110100000100111000001011111000",
   "010000000001001110111000100111010001100000010",
   "010000000001001111010010100111100001100001100",
   "010000000001001111111000100111110001100010110",
   "010000000001010000001010101000000001100100000",
   "010000000001010000111000101000010001100101010",
   "010000000001010001010100101000100001100110100",
   "010000000001010001110010101000110001100111110",
   "010000000001010010011000101001000001101001000",
   "010000000001010010100110101001010001101010011",
   "010000000001010011010110101001100001101011101",
   "010000000001010011101110101001110001101100111",
   "010000000001010100001010101010000001101110010",
   "010000000001010100101010101010010001101111100",
   "010000000001010101001100101010100001110000111",
   "010000000001010101110010101010110001110010010",
   "010000000001010110011010101011000001110011100",
   "010000000001010110101110101011010001110100111",
   "010000000001010111011010101011100001110110010",
   "010000000001010111110000101011110001110111101",
   "010000000001011000011110101100000001111001000",
   "010000000001011000111000101100010001111010011",
   "010000000001011001010110101100100001111011110",
   "010000000001011001101010101100110001111101001",
   "010000000001011010001000101101000001111110100",
   "010000000001011010111110101101010010000000000",
   "010000000001011011011100101101100010000001011",
   "010000000001011011110000101101110010000010111",
   "010000000001011100001110101110000010000100010",
   "010000000001011100101000101110010010000101110",
   "010000000001011101011000101110100010000111001",
   "010000000001011101110100101110110010001000101",
   "010000000001011110000110101111000010001010001",
   "010000000001011110110100101111010010001011100",
   "010000000001011111011110101111100010001101000",
   "010000000001011111110000101111110010001110100",
   "010000000001100000010100110000000010010000000",
   "010000000001100000110100110000010010010001100",
   "010000000001100001010110110000100010010011000",
   "010000000001100001110000110000110010010100100",
   "010000000001100010100010110001000010010110001",
   "010000000001100010101110110001010010010111101",
   "010000000001100011010110110001100010011001001",
   "010000000001100011111100110001110010011010110",
   "010000000001100100010110110010000010011100010",
   "010000000001100100101110110010010010011101111",
   "010000000001100101011010110010100010011111011",
   "010000000001100101111010110010110010100001000",
   "010000000001100110011010110011000010100010101",
   "010000000001100110110010110011010010100100001",
   "010000000001100111011010110011100010100101110",
   "010000000001100111111100110011110010100111011",
   "010000000001101000010100110100000010101001000",
   "010000000001101001000000110100010010101010101",
   "010000000001101001100010110100100010101100010",
   "010000000001101001111010110100110010101110000",
   "010000000001101010001010110101000010101111101",
   "010000000001101010101000110101010010110001010",
   "010000000001101011011100110101100010110010111",
   "010000000001101100000010110101110010110100101",
   "010000000001101100011110110110000010110110010",
   "010000000001101100101110110110010010111000000",
   "010000000001101101001110110110100010111001101",
   "010000000001101101111010110110110010111011011",
   "010000000001101110011010110111000010111101001",
   "010000000001101110110000110111010010111110111",
   "010000000001101111010000110111100011000000100",
   "010000000001110000000000110111110011000010010",
   "010000000001110000100000111000000011000100000",
   "010000000001110000110100111000010011000101110",
   "010000000001110001010100111000100011000111101",
   "010000000001110001111110111000110011001001011",
   "010000000001110010011100111001000011001011001",
   "010000000001110011000100111001010011001100111",
   "010000000001110011010110111001100011001110110",
   "010000000001110011111100111001110011010000100",
   "010000000001110100001000111010000011010010011",
   "010000000001110100111100111010010011010100001",
   "010000000001110101100010111010100011010110000",
   "010000000001110101101110111010110011010111110",
   "010000000001110110001010111011000011011001101",
   "010000000001110110110000111011010011011011100",
   "010000000001110111011000111011100011011101011",
   "010000000001110111101100111011110011011111010",
   "010000000001111000100000111100000011100001001",
   "010000000001111001000010111100010011100011000",
   "010000000001111001010000111100100011100100111",
   "010000000001111010000000111100110011100110110",
   "010000000001111010011000111101000011101000101",
   "010000000001111010110010111101010011101010100",
   "010000000001111011011010111101100011101100100",
   "010000000001111011111110111101110011101110011",
   "010000000001111100001110111110000011110000011",
   "010000000001111100111010111110010011110010010",
   "010000000001111101010000111110100011110100010",
   "010000000001111110000010111110110011110110010",
   "010000000001111110011100111111000011111000001",
   "010000000001111110111000111111010011111010001",
   "010000000001111111010100111111100011111100001",
   "010000000001111111110010111111110011111110001",
   "011111111000000000000000000000000000000000100",
   "000001010000000000000000010000000000000000101",
   "000011100000000000000001000000000000000001111",
   "001000111000000000000010010000000000000101000",
   "010000010000000000000100000000000000001011001",
   "011000100000000000000110010000000000010101011",
   "000011111000000000001001000000000000100100100",
   "010001010000000000001100010000000000111001101",
   "011111100000000000010000000000000001010101111",
   "010000111000000000010100010000000001111010000",
   "000100010000000000011001000000000010100111001",
   "011000101000000000011110010000000011011110011",
   "010000000000000000100100000000000100100000100",
   "001001010000000000101010010000000101101110101",
   "000011101000000000110001000000000111001001111",
   "000001000000000000111000010000001000110011000",
   "011111011000000001000000000000001010101011010",
   "000000110000000001001000010000001100110011011",
   "000100001000000001010001000000001111001100100",
   "001000101000000001011010010000010001110111110",
   "001111111000000001100100000000010100110101111",
   "011000011000000001101110010000011000001000001",
   "000011111000000001111001000000011011101111010",
   "010001010000000010000100010000011111101100011",
   "011111110000000010010000000000100100000000101",
   "010001010000000010011100010000101000101100110",
   "000011110000000010101001000000101101110010000",
   "011001010000000010110110010000110011010001001",
   "001111110000000011000100000000111001001011011",
   "001000011000000011010010010000111111100001101",
   "000100000000000011100001000001000110010100110",
   "000000101000000011110000010001001101100110000",
   "000000010000000100000000000001010101010110001",
   "000000111000000100010000010001011101100110011",
   "000011101000000100100001000001100110010111101",
   "001000100000000100110010010001101111101010111",
   "010000010000000101000100000001111001100001000",
   "011001000000000101010110010010000011111011010",
   "000100000000000101101001000010001110111010100",
   "010000111000000101111100010010011010011111110",
   "011111111000000110010000000010100110101100000",
   "010000111000000110100100010010110011100000010",
   "000100000000000110111001000011000000111101100",
   "011001000000000111001110010011001111000100110",
   "010000010000000111100100000011011101110111000",
   "001001100000000111111010010011101101010101010",
   "000011111000001000010001000011111101100000101",
   "000001001000001000101000010100001110011001111",
   "011111101000001001000000000100100000000010010",
   "000001001000001001011000010100110010011010100",
   "000011110000001001110001000101000101100011111",
   "001001011000001010001010010101011001011111001",
   "010000001000001010100100000101101110001101100",
   "011000111000001010111110010110000011101111111",
   "000011111000001011011001000110011010000111010",
   "010000111000001011110100010110110001010100101",
   "000000000000001100010000000111001001011001000",
   "010001010000001100101100010111100010010101011",
   "000100011000001101001001000111111100001010110",
   "011000111000001101100110011000010110111010010",
   "010000011000001110000100001000110010100100101",
   "001001000000001110100010011001001111001011001",
   "000100110000001111000001001001101100101110100",
   "000001100000001111100000011010001011010000000",
   "000000100000010000000000001010101010110000100",
   "000001101000010000100000011011001011010001000",
   "000100111000010001000001001011101100110010100",
   "001001010000010001100010011100001111010110001",
   "010000110000010010000100001100110010111100101",
   "011001010000010010100110011101010111100111010",
   "000101001000010011001001001101111101010110110",
   "010010000000010011101100011110100100001100011",
   "000001001000010100010000001111001100001001000",
   "010001011000010100110100011111110101001101110",
   "000100110000010101011001010000011111011011011",
   "011001011000010101111110100001001010110011001",
   "010001001000010110100100010001110111010101110",
   "001010001000010111001010100010100101000100100",
   "000101010000010111110001010011010100000000010",
   "000010100000011000011000100100000100001010000",
   "000001000000011001000000010100110101100010111",
   "000001101000011001101000100101101000001011110",
   "000101101000011010010001010110011100000101100",
   "001010101000011010111010100111010001010001011",
   "010001000000011011100100011000000111110000011",
   "011010100000011100001110101000111111100011010",
   "000101010000011100111001011001111000101011010",
   "010010010000011101100100101010110011001001010",
   "000001100000011110010000011011101110111110010",
   "010010111000011110111100101100101100001011010",
   "000101101000011111101001011101101010110001011",
   "011010100000100000010110101110101010110001100",
   "010001110000100001000100011111101100001100101",
   "001011010000100001110010110000101111000011110",
   "000101111000100010100001100001110011011000000",
   "000010111000100011010000110010111001001010010",
   "000010001000100100000000100100000000011011100",
   "000010110000100100110000110101001001001100111",
   "000110100000100101100001100110010011011111001",
   "001011101000100110010010110111011111010011100",
   "010010001000100111000100101000101100101011000",
   "011011110000100111110110111001111011100110011",
   "000110111000101000101001101011001100000110111",
   "010011010000101001011100111100011110001101100",
   "000011000000101010010000101101110001111011000",
   "010100000000101011000100111111000111010000101",
   "000111010000101011111001110000011110001111010",
   "011100000000101100101111000001110110111000000",
   "010011001000101101100100110011010001001011110",
   "001100100000101110011011000100101101001011100",
   "000111011000101111010001110110001010111000011",
   "000100100000110000001001000111101010010011010",
   "000011000000110001000000111001001011011101010",
   "000100111000110001111001001010101110010111001",
   "000111010000110010110001111100010011000010010",
   "001100111000110011101011001101111001011111010",
   "010100000000110100100100111111100001101111011",
   "011100101000110101011111010001001011110011101",
   "000111100000110110011010000010110111101100111",
   "010100111000110111010101010100100101011100001",
   "000100101000111000010001000110010101000010011",
   "010100111000111001001101011000000110100000111",
   "001000101000111010001010001001111001111000010",
   "011101111000111011000111011011101111001001110",
   "010100011000111100000101001101100110010110011",
   "001101100000111101000011011111011111011111000",
   "001001000000111110000010010001011010100100101",
   "000110001000111111000001100011010111101000011",
   "000100101001000000000001010101010110101011010",
   "000110101001000001000001100111010111101110000",
   "001001010001000010000010011001011010110010000",
   "001110011001000011000011101011011111111000000",
   "010101111001000100000101011101100111000001000",
   "011111000001000101000111101111110000001110001",
   "001001110001000110001010100001111011100000011",
   "010111000001000111001101110100001000111000101",
   "000101110001001000010001100110011000011000000",
   "010111001001001001010101111000101001111111011",
   "001010000001001010011010101010111101101111111",
   "011111101001001011011111111101010011101010011",
   "010110101001001100100101101111101011110000000",
   "010000011001001101101100000010000110000001101",
   "001010101001001110110010110100100010100000100",
   "001000101001001111111010000111000001001101010",
   "000111010001010001000001111001100010001001010",
   "001000011001010010001010001100000101010101010",
   "001100001001010011010010111110101010110010010",
   "010000110001010100011100010001010010100001100",
   "010111111001010101100110000011111100100011110",
   "000001110001010110110000010110101000111010000",
   "001100010001010111111011001001010111100101100",
   "011001011001011001000110011100001000100111000",
   "001000010001011010010010001110111011111111101",
   "011001111001011011011110100001110001110000010",
   "001101010001011100101011010100101001111010000",
   "000010010001011101111000100111100100011101111",
   "011001000001011111000110011010100001011100111",
   "010010100001100000010100101101100000110111111",
   "001101111001100001100011100000100010110000000",
   "001010111001100010110010110011100111000110010",
   "001010101001100100000010100110101101111011100",
   "001011010001100101010010111001110111010001000",
   "001110101001100110100011101101000011000111100",
   "010011111001100111110101000000010001100000001",
   "011010111001101001000110110011100010011011111",
   "000100110001101010011001000110110101111011101",
   "001111011001101011101011111010001100000000101",
   "011100111001101100111111001101100100101011101",
   "001100010001101110010011000000111111111101110",
   "011101100001101111100111010100011101111000000",
   "010000101001110000111100000111111110011011011",
   "000101101001110010010001011011100001101000111",
   "011100100001110011100111001111000111100001100",
   "010110010001110100111101100010110000000110001",
   "010001000001110110010100010110011011011000000",
   "001110101001110111101011101010001001010111111",
   "001101010001111001000011011101111010000111000",
   "001110110001111010011011110001101101100110001",
   "010010001001111011110100100101100011110110011",
   "010111110001111101001101111001011100111000110",
   "011111001001111110100111101101011000101110010",
   "000111100010000000000010000001010111011000000",
   "010010111010000001011100110101011000110110110",
   "000000100010000010111000001001011101001011101",
   "001111111010000100010011111101100100010111101",
   "000001011010000101110000010001101110011011110",
   "010100000010000111001101000101111011011001001",
   "001001100010001000101010011010001011010000100",
   "000001010010001010001000001110011110000011000",
   "011010000010001011100110100010110011110001110",
   "010100111010001101000101010111001100011101101",
   "010010110010001110100100101011101000000111100",
   "010001111010010000000100100000000110110000101",
   "010011001010010001100100110100101000011001111",
   "010110011010010011000101101001001101000100010",
   "011011111010010100100110111101110100110000110",
   "000010100010010110001000110010011111100000100",
   "001100100010010111101011000111001101010100010",
   "010111100010011001001101111011111110001101010",
   "000100101010011010110001010000110010001100011",
   "010100001010011100010101000101101001010010101",
   "000101110010011101111001011010100011100001000",
   "011000101010011111011110001111100000111000101",
   "001101111010100001000011100100100001011010011",
   "000101010010100010101001011001100101000111010",
   "011110111010100100001111101110101100000000010",
   "011001111010100101110110100011110110000110100",
   "010111001010100111011101111001000011011010111",
   "010110110010101001000101101110010011111110011",
   "010111101010101010101110000011100111110010001",
   "011010111010101100010110111000111110110111000",
   "000000100010101110000000001110011001001110000",
   "001000100010101111101010000011110110111000001",
   "010001111010110001010100011001010111110110100",
   "011100100010110010111111001110111100001010001",
   "001001101010110100101010100100100011110011111",
   "011001001010110110010110011010001110110100110",
   "001011001010111000000010101111111101001101110",
   "011110100010111001101111100101101111000000000",
   "010011011010111011011100111011100100001100100",
   "001010110010111101001010110001011100110100001",
   "000100100010111110111001000111011000110111111",
   "011111111011000000100111111101011000011000111",
   "011100101011000010010111010011011011011000001",
   "011100000011000100000111001001100001110110100",
   "011101111011000101110111011111101011110101000",
   "000001010011000111101000010101111001010100110",
   "000110010011001001011001101100001010010110110",
   "001101110011001011001011100010011110111011111",
   "010110111011001100111101111000110111000101010",
   "000010110011001110110000101111010010110011110",
   "010000000011010000100100000101110010001000100",
   "000000001011010010010111111100010101000100011",
   "010000110011010100001100010010111011101000101",
   "000100000011010110000001001001100101110110000",
   "011010001011010111110110100000010011101101100",
   "010001110011011001101100010111000101010000010",
   "001011000011011011100010101101111010011111010",
   "000110001011011101011001100100110011011011100",
   "000100000011011111010000111011110000000101111",
   "000010101011100001001000110010110000011111101",
   "000100000011100011000001001001110100101001100",
   "001000001011100100111010000000111100100100100",
   "001101000011100110110011011000001000010001111",
   "010100110011101000101101001111010111110010011",
   "011110011011101010100111100110101011000111001",
   "001001101011101100100010011110000010010001001",
   "010110111011101110011101110101011101010001011",
   "000111000011110000011001101100111100001000110",
   "011000000011110010010110000100011110111000100",
   "001011111011110100010010111100000101100001011",
   "000000101011110110010000010011110000000100101",
   "011000011011111000001110001011011110100011000",
   "010010000011111010001100100011010000111101101",
   "001101101011111100001011011011000111010101100",
   "001011010011111110001010110011000001101011101",
      others => (others => '0'));
      	begin 
      return tmp;
      end init_rom;
	signal rom : memory_t := init_rom;
   signal Y1 :  std_logic_vector(44 downto 0);
   signal Y0 :  std_logic_vector(44 downto 0);
   signal Z1 :  std_logic_vector(8 downto 0);
   signal Z0 :  std_logic_vector(8 downto 0);
begin
Z0 <= '1' & X;
Z1 <= '0' & X;
	process(clk)
   begin
   if(rising_edge(clk)) then
     if(Enable='1') then
   	Y1 <= rom(  TO_INTEGER(unsigned(Z1)));
   	Y0 <= rom(  TO_INTEGER(unsigned(Z0)));
     end if;
   end if;
   end process;
    Y <= Y1 & Y0(43 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                            FunctionEvaluator_68
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Mioara Joldes, Florent de Dinechin (2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FunctionEvaluator_68 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(32 downto 0);
          R_old : out  std_logic_vector(33 downto 0);
          R : out  std_logic_vector(33 downto 0)   );
end entity;

architecture arch of FunctionEvaluator_68 is
   component PolyCoeffTable_8_89 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             X : in  std_logic_vector(7 downto 0);
             Y : out  std_logic_vector(88 downto 0)   );
   end component;

   component PolynomialEvaluator_degree2_uid71 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             Y : in  std_logic_vector(24 downto 0);
             a0 : in  std_logic_vector(35 downto 0);
             a1 : in  std_logic_vector(29 downto 0);
             a2 : in  std_logic_vector(22 downto 0);
             R_old : out  std_logic_vector(36 downto 0);
             R : out  std_logic_vector(36 downto 0)   );
   end component;

signal addr :  std_logic_vector(7 downto 0);
signal Coef, Coef_d1 :  std_logic_vector(88 downto 0);
signal y :  std_logic_vector(24 downto 0);
signal a0 :  std_logic_vector(35 downto 0);
signal a1 :  std_logic_vector(29 downto 0);
signal a2 :  std_logic_vector(22 downto 0);
signal Rpe :  std_logic_vector(36 downto 0);
signal Rpe_old :  std_logic_vector(36 downto 0);

signal X_d1, X_d2 :  std_logic_vector(32 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
           if(Enable='1') then
            Coef_d1 <=  Coef;
            X_d1 <=  X;
            X_d2 <=  X_d1;
           end if;
         end if;
      end process;
   addr <= X(32 downto 25);
   GeneratedTable: PolyCoeffTable_8_89  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 X => addr,
                 Y => Coef);
   ----------------Synchro barrier, entering cycle 1----------------
   ----------------Synchro barrier, entering cycle 2----------------
   y <= X_d2(24 downto 0);
   a0<= Coef_d1(35 downto 0);
   a1<= Coef_d1(65 downto 36);
   a2<= Coef_d1(88 downto 66);
   PolynomialEvaluator: PolynomialEvaluator_degree2_uid71  -- pipelineDepth=8 maxInDelay=0
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 R => Rpe,
                 R_old => Rpe_old,
                 Y => y,
                 a0 => a0,
                 a1 => a1,
                 a2 => a2);
   ----------------Synchro barrier, entering cycle 10----------------
   -- weight of poly result is : 1
    R_old <= Rpe_old(36 downto 3);
    R <= Rpe(36 downto 3);
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_12_f400_uid40
--                     (IntAdderClassical_12_f400_uid42)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_12_f400_uid40 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL     rst : in std_logic;
          X : in  std_logic_vector(11 downto 0);
          Y : in  std_logic_vector(11 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of IntAdder_12_f400_uid40 is
signal X_d1 :  std_logic_vector(11 downto 0);
signal Y_d1 :  std_logic_vector(11 downto 0);
signal Cin_d1 : std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
           if(Enable='1') then
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
           end if;
         end if;
      end process;
   --Classical
   ----------------Synchro barrier, entering cycle 1----------------
    R <= X_d1 + Y_d1 + Cin_d1;
end architecture;
--------------------------------------------------------------------------------
--                 FixRealKCM_M3_6_0_1_log_2_unsigned_Table_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity FixRealKCM_M3_6_0_1_log_2_unsigned_Table_1 is
   port (-- OL clk, rst : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of FixRealKCM_M3_6_0_1_log_2_unsigned_Table_1 is
begin
  with X select  Y <= 
   "000000001000" when "0000",
   "000011000001" when "0001",
   "000101111001" when "0010",
   "001000110010" when "0011",
   "001011101011" when "0100",
   "001110100011" when "0101",
   "010001011100" when "0110",
   "010100010101" when "0111",
   "010111001101" when "1000",
   "011010000110" when "1001",
   "011100111111" when "1010",
   "011111110111" when "1011",
   "100010110000" when "1100",
   "100101101001" when "1101",
   "101000100001" when "1110",
   "101011011010" when "1111",
   "------------" when others;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_M3_6_0_1_log_2_unsigned_Table_0
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity FixRealKCM_M3_6_0_1_log_2_unsigned_Table_0 is
   port (-- OL clk, rst : in std_logic;
          X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(7 downto 0)   );
end entity;

architecture arch of FixRealKCM_M3_6_0_1_log_2_unsigned_Table_0 is
begin
  with X select  Y <= 
   "00000000" when "000000",
   "00000011" when "000001",
   "00000110" when "000010",
   "00001001" when "000011",
   "00001100" when "000100",
   "00001110" when "000101",
   "00010001" when "000110",
   "00010100" when "000111",
   "00010111" when "001000",
   "00011010" when "001001",
   "00011101" when "001010",
   "00100000" when "001011",
   "00100011" when "001100",
   "00100110" when "001101",
   "00101000" when "001110",
   "00101011" when "001111",
   "00101110" when "010000",
   "00110001" when "010001",
   "00110100" when "010010",
   "00110111" when "010011",
   "00111010" when "010100",
   "00111101" when "010101",
   "00111111" when "010110",
   "01000010" when "010111",
   "01000101" when "011000",
   "01001000" when "011001",
   "01001011" when "011010",
   "01001110" when "011011",
   "01010001" when "011100",
   "01010100" when "011101",
   "01010111" when "011110",
   "01011001" when "011111",
   "01011100" when "100000",
   "01011111" when "100001",
   "01100010" when "100010",
   "01100101" when "100011",
   "01101000" when "100100",
   "01101011" when "100101",
   "01101110" when "100110",
   "01110001" when "100111",
   "01110011" when "101000",
   "01110110" when "101001",
   "01111001" when "101010",
   "01111100" when "101011",
   "01111111" when "101100",
   "10000010" when "101101",
   "10000101" when "101110",
   "10001000" when "101111",
   "10001010" when "110000",
   "10001101" when "110001",
   "10010000" when "110010",
   "10010011" when "110011",
   "10010110" when "110100",
   "10011001" when "110101",
   "10011100" when "110110",
   "10011111" when "110111",
   "10100010" when "111000",
   "10100100" when "111001",
   "10100111" when "111010",
   "10101010" when "111011",
   "10101101" when "111100",
   "10110000" when "111101",
   "10110011" when "111110",
   "10110110" when "111111",
   "--------" when others;
end architecture;

--------------------------------------------------------------------------------
--                     FixRealKCM_M3_6_0_1_log_2_unsigned
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_M3_6_0_1_log_2_unsigned is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL     rst : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          R : out  std_logic_vector(7 downto 0)   );
end entity;

architecture arch of FixRealKCM_M3_6_0_1_log_2_unsigned is
   component FixRealKCM_M3_6_0_1_log_2_unsigned_Table_0 is
      port ( -- OL clk, rst : in std_logic;
             X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(7 downto 0)   );
   end component;

   component FixRealKCM_M3_6_0_1_log_2_unsigned_Table_1 is
      port (-- OL  clk, rst : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(11 downto 0)   );
   end component;

   component IntAdder_12_f400_uid40 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL        rst : in std_logic;
             X : in  std_logic_vector(11 downto 0);
             Y : in  std_logic_vector(11 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(11 downto 0)   );
   end component;

signal d0 :  std_logic_vector(5 downto 0);
signal pp0 :  std_logic_vector(7 downto 0);
signal addOp0 :  std_logic_vector(11 downto 0);
signal d1 :  std_logic_vector(3 downto 0);
signal pp1 :  std_logic_vector(11 downto 0);
signal addOp1 :  std_logic_vector(11 downto 0);
signal OutRes :  std_logic_vector(11 downto 0);
constant zero : std_logic := '0';
attribute rom_extract: string;
attribute rom_style: string;
attribute rom_extract of FixRealKCM_M3_6_0_1_log_2_unsigned_Table_0: component is "yes";
attribute rom_extract of FixRealKCM_M3_6_0_1_log_2_unsigned_Table_1: component is "yes";
attribute rom_style of FixRealKCM_M3_6_0_1_log_2_unsigned_Table_0: component is "distributed";
attribute rom_style of FixRealKCM_M3_6_0_1_log_2_unsigned_Table_1: component is "distributed";
begin
--   process(clk)
--      begin
--         if clk'event and clk = '1' then
--         end if;
--      end process;
   d0 <= X(5 downto 0);
   KCMTable_0: FixRealKCM_M3_6_0_1_log_2_unsigned_Table_0  -- pipelineDepth=0 maxInDelay=0
      port map (-- OL  clk  => clk,
                -- OL rst  => rst,
                 X => d0,
                 Y => pp0);
   addOp0 <= (11 downto 8 => '0') & pp0;
   d1 <= X(9 downto 6);
   KCMTable_1: FixRealKCM_M3_6_0_1_log_2_unsigned_Table_1  -- pipelineDepth=0 maxInDelay=0
      port map (-- OL clk  => clk,
                -- OL rst  => rst,
                 X => d1,
                 Y => pp1);
   addOp1 <= pp1;
   Result_Adder: IntAdder_12_f400_uid40  -- pipelineDepth=1 maxInDelay=1.80264e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 Cin => zero,
                 R => OutRes,
                 X => addOp0,
                 Y => addOp1);
   ----------------Synchro barrier, entering cycle 1----------------
   R <= OutRes(11 downto 4);
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_59_f400_uid55
--                     (IntAdderClassical_59_f400_uid57)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_59_f400_uid55 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(58 downto 0);
          Y : in  std_logic_vector(58 downto 0);
          Cin : in std_logic;
          R : out  std_logic_vector(58 downto 0)   );
end entity;

architecture arch of IntAdder_59_f400_uid55 is
signal x0 :  std_logic_vector(41 downto 0);
signal y0 :  std_logic_vector(41 downto 0);
signal x1, x1_d1 :  std_logic_vector(16 downto 0);
signal y1, y1_d1 :  std_logic_vector(16 downto 0);
signal sum0, sum0_d1 :  std_logic_vector(42 downto 0);
signal sum1 :  std_logic_vector(17 downto 0);
signal X_d1 :  std_logic_vector(58 downto 0);
signal Y_d1 :  std_logic_vector(58 downto 0);
signal Cin_d1 : std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
           if(Enable='1') then
            x1_d1 <=  x1;
            y1_d1 <=  y1;
            sum0_d1 <=  sum0;
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
           end if;
         end if;
      end process;
   --Classical
   ----------------Synchro barrier, entering cycle 1----------------
   x0 <= X_d1(41 downto 0);
   y0 <= Y_d1(41 downto 0);
   x1 <= X_d1(58 downto 42);
   y1 <= Y_d1(58 downto 42);
   sum0 <= ( "0" & x0) + ( "0" & y0)  + Cin_d1;
   ----------------Synchro barrier, entering cycle 2----------------
   sum1 <= ( "0" & x1_d1) + ( "0" & y1_d1)  + sum0_d1(42);
   R <= sum1(16 downto 0) & sum0_d1(41 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_0_7_M51_log_2_unsigned_Table_1
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity FixRealKCM_0_7_M51_log_2_unsigned_Table_1 is
   port (-- OL clk, rst : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : out  std_logic_vector(58 downto 0)   );
end entity;

architecture arch of FixRealKCM_0_7_M51_log_2_unsigned_Table_1 is
begin
  with X select  Y <= 
   "00000000000000000000000000000000000000000000000000000000000" when "00",
   "00101100010111001000010111111101111101000111001111011110011" when "01",
   "01011000101110010000101111111011111010001110011110111100111" when "10",
   "10000101000101011001000111111001110111010101101110011011010" when "11",
   "-----------------------------------------------------------" when others;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_0_7_M51_log_2_unsigned_Table_0
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
entity FixRealKCM_0_7_M51_log_2_unsigned_Table_0 is
   port (
-- OL clk, rst : in std_logic;
          X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(56 downto 0)   );
end entity;

architecture arch of FixRealKCM_0_7_M51_log_2_unsigned_Table_0 is
begin
  with X select  Y <= 
   "000000000000000000000000000000000000000000000000000000000" when "000000",
   "000000101100010111001000010111111101111101000111001111100" when "000001",
   "000001011000101110010000101111111011111010001110011111000" when "000010",
   "000010000101000101011001000111111001110111010101101110011" when "000011",
   "000010110001011100100001011111110111110100011100111101111" when "000100",
   "000011011101110011101001110111110101110001100100001101011" when "000101",
   "000100001010001010110010001111110011101110101011011100111" when "000110",
   "000100110110100001111010100111110001101011110010101100011" when "000111",
   "000101100010111001000010111111101111101000111001111011110" when "001000",
   "000110001111010000001011010111101101100110000001001011010" when "001001",
   "000110111011100111010011101111101011100011001000011010110" when "001010",
   "000111100111111110011100000111101001100000001111101010010" when "001011",
   "001000010100010101100100011111100111011101010110111001110" when "001100",
   "001001000000101100101100110111100101011010011110001001001" when "001101",
   "001001101101000011110101001111100011010111100101011000101" when "001110",
   "001010011001011010111101100111100001010100101100101000001" when "001111",
   "001011000101110010000101111111011111010001110011110111101" when "010000",
   "001011110010001001001110010111011101001110111011000111001" when "010001",
   "001100011110100000010110101111011011001100000010010110100" when "010010",
   "001101001010110111011111000111011001001001001001100110000" when "010011",
   "001101110111001110100111011111010111000110010000110101100" when "010100",
   "001110100011100101101111110111010101000011011000000101000" when "010101",
   "001111001111111100111000001111010011000000011111010100100" when "010110",
   "001111111100010100000000100111010000111101100110100011111" when "010111",
   "010000101000101011001000111111001110111010101101110011011" when "011000",
   "010001010101000010010001010111001100110111110101000010111" when "011001",
   "010010000001011001011001101111001010110100111100010010011" when "011010",
   "010010101101110000100010000111001000110010000011100001111" when "011011",
   "010011011010000111101010011111000110101111001010110001010" when "011100",
   "010100000110011110110010110111000100101100010010000000110" when "011101",
   "010100110010110101111011001111000010101001011001010000010" when "011110",
   "010101011111001101000011100111000000100110100000011111110" when "011111",
   "010110001011100100001011111110111110100011100111101111010" when "100000",
   "010110110111111011010100010110111100100000101110111110101" when "100001",
   "010111100100010010011100101110111010011101110110001110001" when "100010",
   "011000010000101001100101000110111000011010111101011101101" when "100011",
   "011000111101000000101101011110110110011000000100101101001" when "100100",
   "011001101001010111110101110110110100010101001011111100101" when "100101",
   "011010010101101110111110001110110010010010010011001100000" when "100110",
   "011011000010000110000110100110110000001111011010011011100" when "100111",
   "011011101110011101001110111110101110001100100001101011000" when "101000",
   "011100011010110100010111010110101100001001101000111010100" when "101001",
   "011101000111001011011111101110101010000110110000001010000" when "101010",
   "011101110011100010101000000110101000000011110111011001011" when "101011",
   "011110011111111001110000011110100110000000111110101000111" when "101100",
   "011111001100010000111000110110100011111110000101111000011" when "101101",
   "011111111000101000000001001110100001111011001101000111111" when "101110",
   "100000100100111111001001100110011111111000010100010111011" when "101111",
   "100001010001010110010001111110011101110101011011100110111" when "110000",
   "100001111101101101011010010110011011110010100010110110010" when "110001",
   "100010101010000100100010101110011001101111101010000101110" when "110010",
   "100011010110011011101011000110010111101100110001010101010" when "110011",
   "100100000010110010110011011110010101101001111000100100110" when "110100",
   "100100101111001001111011110110010011100110111111110100010" when "110101",
   "100101011011100001000100001110010001100100000111000011101" when "110110",
   "100110000111111000001100100110001111100001001110010011001" when "110111",
   "100110110100001111010100111110001101011110010101100010101" when "111000",
   "100111100000100110011101010110001011011011011100110010001" when "111001",
   "101000001100111101100101101110001001011000100100000001101" when "111010",
   "101000111001010100101110000110000111010101101011010001000" when "111011",
   "101001100101101011110110011110000101010010110010100000100" when "111100",
   "101010010010000010111110110110000011001111111001110000000" when "111101",
   "101010111110011010000111001110000001001101000000111111100" when "111110",
   "101011101010110001001111100101111111001010001000001111000" when "111111",
   "---------------------------------------------------------" when others;
end architecture;

--------------------------------------------------------------------------------
--                     FixRealKCM_0_7_M51_log_2_unsigned
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_0_7_M51_log_2_unsigned is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL, rst : in std_logic;
          X : in  std_logic_vector(7 downto 0);
          R : out  std_logic_vector(58 downto 0)   );
end entity;

architecture arch of FixRealKCM_0_7_M51_log_2_unsigned is
   component FixRealKCM_0_7_M51_log_2_unsigned_Table_0 is
      port ( -- OL clk : in std_logic;
             -- OL Enable : in std_logic;
-- OL, rst : in std_logic;
             X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(56 downto 0)   );
   end component;

   component FixRealKCM_0_7_M51_log_2_unsigned_Table_1 is
      port (
-- OL clk : in std_logic;
-- OL             Enable : in std_logic;
-- OL, rst : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : out  std_logic_vector(58 downto 0)   );
   end component;

   component IntAdder_59_f400_uid55 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL , rst : in std_logic;
             X : in  std_logic_vector(58 downto 0);
             Y : in  std_logic_vector(58 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(58 downto 0)   );
   end component;

signal d0 :  std_logic_vector(5 downto 0);
signal pp0 :  std_logic_vector(56 downto 0);
signal addOp0 :  std_logic_vector(58 downto 0);
signal d1 :  std_logic_vector(1 downto 0);
signal pp1 :  std_logic_vector(58 downto 0);
signal addOp1 :  std_logic_vector(58 downto 0);
signal OutRes :  std_logic_vector(58 downto 0);
attribute rom_extract: string;
attribute rom_style: string;
attribute rom_extract of FixRealKCM_0_7_M51_log_2_unsigned_Table_0: component is "yes";
attribute rom_extract of FixRealKCM_0_7_M51_log_2_unsigned_Table_1: component is "yes";
attribute rom_style of FixRealKCM_0_7_M51_log_2_unsigned_Table_0: component is "distributed";
attribute rom_style of FixRealKCM_0_7_M51_log_2_unsigned_Table_1: component is "distributed";
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   d0 <= X(5 downto 0);
   KCMTable_0: FixRealKCM_0_7_M51_log_2_unsigned_Table_0  -- pipelineDepth=0 maxInDelay=0
      port map (
-- OL clk  => clk,
-- OL                 Enable => Enable,
-- OL                 rst  => rst,
                 X => d0,
                 Y => pp0);
   addOp0 <= (58 downto 57 => '0') & pp0;
   d1 <= X(7 downto 6);
   KCMTable_1: FixRealKCM_0_7_M51_log_2_unsigned_Table_1  -- pipelineDepth=0 maxInDelay=0
      port map (-- OL clk  => clk,
-- OL                 Enable => Enable,
-- OL                 rst  => rst,
                 X => d1,
                 Y => pp1);
   addOp1 <= pp1;
   Result_Adder: IntAdder_59_f400_uid55  -- pipelineDepth=2 maxInDelay=2.35544e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 Cin => '0',
                 R => OutRes,
                 X => addOp0,
                 Y => addOp1);
   ----------------Synchro barrier, entering cycle 2----------------
   R <= OutRes(58 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                               FPExp_8_47_400
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, Bogdan Pasca (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 32 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPExp_8_47_400 is
   port ( clk : in std_logic;
          Enable : in std_logic;
-- OL , rst : in std_logic;
          X : in  std_logic_vector(8+47+2 downto 0);
          R : out  std_logic_vector(8+47+2 downto 0)   );
end entity;

architecture arch of FPExp_8_47_400 is
   component FixRealKCM_0_7_M51_log_2_unsigned is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             X : in  std_logic_vector(7 downto 0);
             R : out  std_logic_vector(58 downto 0)   );
   end component;

   component FixRealKCM_M3_6_0_1_log_2_unsigned is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             R : out  std_logic_vector(7 downto 0)   );
   end component;

   component FunctionEvaluator_68 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             X : in  std_logic_vector(32 downto 0);
             R_old : out  std_logic_vector(33 downto 0);
             R : out  std_logic_vector(33 downto 0)   );
   end component;

   component IntAdder_43_f400_uid107 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             X : in  std_logic_vector(42 downto 0);
             Y : in  std_logic_vector(42 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(42 downto 0)   );
   end component;

   component IntAdder_43_f400_uid113 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             X : in  std_logic_vector(42 downto 0);
             Y : in  std_logic_vector(42 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(42 downto 0)   );
   end component;

   component IntAdder_51_f484_uid61 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             X : in  std_logic_vector(50 downto 0);
             Y : in  std_logic_vector(50 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(50 downto 0)   );
   end component;

   component IntAdder_52_f400_uid133 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             X : in  std_logic_vector(51 downto 0);
             Y : in  std_logic_vector(51 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(51 downto 0)   );
   end component;

   component IntAdder_57_f400_uid139 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL , rst : in std_logic;
             X : in  std_logic_vector(56 downto 0);
             Y : in  std_logic_vector(56 downto 0);
             Cin : in std_logic;
             R : out  std_logic_vector(56 downto 0)   );
   end component;

   component IntMultiplier_42_43_unsigned_uid119 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             X : in  std_logic_vector(41 downto 0);
             Y : in  std_logic_vector(42 downto 0);
             R : out  std_logic_vector(84 downto 0)   );
   end component;

   component LeftShifter_48_by_max_58_uid41 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL, rst : in std_logic;
             X : in  std_logic_vector(47 downto 0);
             S : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(105 downto 0)   );
   end component;

   component firstExpTable_9_52 is
      port ( clk : in std_logic;
             Enable : in std_logic;
-- OL , rst : in std_logic;
             X : in  std_logic_vector(8 downto 0);
             Y : out  std_logic_vector(51 downto 0)   );
   end component;

signal Xexn, Xexn_d1, Xexn_d2, Xexn_d3, Xexn_d4, Xexn_d5, Xexn_d6, Xexn_d7, Xexn_d8, Xexn_d9, Xexn_d10, Xexn_d11, Xexn_d12, Xexn_d13, Xexn_d14, Xexn_d15, Xexn_d16, Xexn_d17, Xexn_d18, Xexn_d19, Xexn_d20, Xexn_d21, Xexn_d22, Xexn_d23, Xexn_d24, Xexn_d25, Xexn_d26, Xexn_d27, Xexn_d28, Xexn_d29, Xexn_d30, Xexn_d31, Xexn_d32 :  std_logic_vector(1 downto 0);
signal XSign, XSign_d1, XSign_d2, XSign_d3, XSign_d4, XSign_d5, XSign_d6, XSign_d7, XSign_d8, XSign_d9, XSign_d10, XSign_d11, XSign_d12, XSign_d13, XSign_d14, XSign_d15, XSign_d16, XSign_d17, XSign_d18, XSign_d19, XSign_d20, XSign_d21, XSign_d22, XSign_d23, XSign_d24, XSign_d25, XSign_d26, XSign_d27, XSign_d28, XSign_d29, XSign_d30, XSign_d31, XSign_d32 : std_logic;
signal XexpField :  std_logic_vector(7 downto 0);
signal Xfrac :  std_logic_vector(46 downto 0);
signal e0 :  std_logic_vector(9 downto 0);
signal shiftVal, shiftVal_d1 :  std_logic_vector(9 downto 0);
signal resultWillBeOne, resultWillBeOne_d1, resultWillBeOne_d2, resultWillBeOne_d3 : std_logic;
signal mXu :  std_logic_vector(47 downto 0);
signal oufl0, oufl0_d1, oufl0_d2, oufl0_d3, oufl0_d4, oufl0_d5, oufl0_d6, oufl0_d7, oufl0_d8, oufl0_d9, oufl0_d10, oufl0_d11, oufl0_d12, oufl0_d13, oufl0_d14, oufl0_d15, oufl0_d16, oufl0_d17, oufl0_d18, oufl0_d19, oufl0_d20, oufl0_d21, oufl0_d22, oufl0_d23, oufl0_d24, oufl0_d25, oufl0_d26, oufl0_d27, oufl0_d28, oufl0_d29, oufl0_d30, oufl0_d31 : std_logic;
signal shiftValIn :  std_logic_vector(5 downto 0);
signal fixX0, fixX0_d1 :  std_logic_vector(105 downto 0);
signal fixX, fixX_d1, fixX_d2, fixX_d3 :  std_logic_vector(58 downto 0);
signal xMulIn :  std_logic_vector(9 downto 0);
signal absK, absK_d1 :  std_logic_vector(7 downto 0);
signal minusAbsK :  std_logic_vector(8 downto 0);
signal K, K_d1, K_d2, K_d3, K_d4, K_d5, K_d6, K_d7, K_d8, K_d9, K_d10, K_d11, K_d12, K_d13, K_d14, K_d15, K_d16, K_d17, K_d18, K_d19, K_d20, K_d21, K_d22, K_d23, K_d24, K_d25 :  std_logic_vector(8 downto 0);
signal absKLog2 :  std_logic_vector(58 downto 0);
signal subOp1 :  std_logic_vector(50 downto 0);
signal subOp2 :  std_logic_vector(50 downto 0);
signal Y :  std_logic_vector(50 downto 0);
signal Addr1 :  std_logic_vector(8 downto 0);
signal Z, Z_d1, Z_d2, Z_d3, Z_d4, Z_d5, Z_d6, Z_d7, Z_d8, Z_d9, Z_d10, Z_d11 :  std_logic_vector(41 downto 0);
signal Zhigh, Zhigh_d1 :  std_logic_vector(32 downto 0);
signal expA, expA_d1, expA_d2, expA_d3, expA_d4, expA_d5, expA_d6, expA_d7, expA_d8, expA_d9, expA_d10, expA_d11, expA_d12, expA_d13, expA_d14, expA_d15, expA_d16, expA_d17, expA_d18 :  std_logic_vector(51 downto 0);
signal expZmZm1_0 :  std_logic_vector(33 downto 0);
signal expZmZm1 :  std_logic_vector(33 downto 0);
signal expZminus1X :  std_logic_vector(42 downto 0);
signal expZminus1Y :  std_logic_vector(42 downto 0);
signal expZminus1 :  std_logic_vector(42 downto 0);
signal expArounded0 :  std_logic_vector(42 downto 0);
signal expArounded, expArounded_d1, expArounded_d2, expArounded_d3, expArounded_d4, expArounded_d5, expArounded_d6, expArounded_d7, expArounded_d8, expArounded_d9, expArounded_d10 :  std_logic_vector(41 downto 0);
signal lowerProduct :  std_logic_vector(84 downto 0);
signal extendedLowerProduct :  std_logic_vector(51 downto 0);
signal expY :  std_logic_vector(51 downto 0);
signal needNoNorm : std_logic;
signal preRoundBiasSig :  std_logic_vector(56 downto 0);
signal roundBit : std_logic;
signal roundNormAddend :  std_logic_vector(56 downto 0);
signal roundedExpSigRes :  std_logic_vector(56 downto 0);
signal roundedExpSig :  std_logic_vector(56 downto 0);
signal ofl1 : std_logic;
signal ofl2 : std_logic;
signal ofl3 : std_logic;
signal ofl : std_logic;
signal ufl1 : std_logic;
signal ufl2 : std_logic;
signal ufl3 : std_logic;
signal ufl : std_logic;
signal Rexn :  std_logic_vector(1 downto 0);
constant g: positive := 4;
constant wE: positive := 8;
constant wF: positive := 47;
constant wFIn: positive := 47;

signal  expZmZm1_0_old :  std_logic_vector(33 downto 0);

signal Tmp :  std_logic_vector(58 downto 0);

begin
   process(clk)
      begin
         if clk'event and clk = '1' then
           if(Enable='1') then
            Xexn_d1 <=  Xexn;
            Xexn_d2 <=  Xexn_d1;
            Xexn_d3 <=  Xexn_d2;
            Xexn_d4 <=  Xexn_d3;
            Xexn_d5 <=  Xexn_d4;
            Xexn_d6 <=  Xexn_d5;
            Xexn_d7 <=  Xexn_d6;
            Xexn_d8 <=  Xexn_d7;
            Xexn_d9 <=  Xexn_d8;
            Xexn_d10 <=  Xexn_d9;
            Xexn_d11 <=  Xexn_d10;
            Xexn_d12 <=  Xexn_d11;
            Xexn_d13 <=  Xexn_d12;
            Xexn_d14 <=  Xexn_d13;
            Xexn_d15 <=  Xexn_d14;
            Xexn_d16 <=  Xexn_d15;
            Xexn_d17 <=  Xexn_d16;
            Xexn_d18 <=  Xexn_d17;
            Xexn_d19 <=  Xexn_d18;
            Xexn_d20 <=  Xexn_d19;
            Xexn_d21 <=  Xexn_d20;
            Xexn_d22 <=  Xexn_d21;
            Xexn_d23 <=  Xexn_d22;
            Xexn_d24 <=  Xexn_d23;
            Xexn_d25 <=  Xexn_d24;
            Xexn_d26 <=  Xexn_d25;
            Xexn_d27 <=  Xexn_d26;
            Xexn_d28 <=  Xexn_d27;
            Xexn_d29 <=  Xexn_d28;
            Xexn_d30 <=  Xexn_d29;
            Xexn_d31 <=  Xexn_d30;
            Xexn_d32 <=  Xexn_d31;
            XSign_d1 <=  XSign;
            XSign_d2 <=  XSign_d1;
            XSign_d3 <=  XSign_d2;
            XSign_d4 <=  XSign_d3;
            XSign_d5 <=  XSign_d4;
            XSign_d6 <=  XSign_d5;
            XSign_d7 <=  XSign_d6;
            XSign_d8 <=  XSign_d7;
            XSign_d9 <=  XSign_d8;
            XSign_d10 <=  XSign_d9;
            XSign_d11 <=  XSign_d10;
            XSign_d12 <=  XSign_d11;
            XSign_d13 <=  XSign_d12;
            XSign_d14 <=  XSign_d13;
            XSign_d15 <=  XSign_d14;
            XSign_d16 <=  XSign_d15;
            XSign_d17 <=  XSign_d16;
            XSign_d18 <=  XSign_d17;
            XSign_d19 <=  XSign_d18;
            XSign_d20 <=  XSign_d19;
            XSign_d21 <=  XSign_d20;
            XSign_d22 <=  XSign_d21;
            XSign_d23 <=  XSign_d22;
            XSign_d24 <=  XSign_d23;
            XSign_d25 <=  XSign_d24;
            XSign_d26 <=  XSign_d25;
            XSign_d27 <=  XSign_d26;
            XSign_d28 <=  XSign_d27;
            XSign_d29 <=  XSign_d28;
            XSign_d30 <=  XSign_d29;
            XSign_d31 <=  XSign_d30;
            XSign_d32 <=  XSign_d31;
            shiftVal_d1 <=  shiftVal;
            resultWillBeOne_d1 <=  resultWillBeOne;
            resultWillBeOne_d2 <=  resultWillBeOne_d1;
            resultWillBeOne_d3 <=  resultWillBeOne_d2;
            oufl0_d1 <=  oufl0;
            oufl0_d2 <=  oufl0_d1;
            oufl0_d3 <=  oufl0_d2;
            oufl0_d4 <=  oufl0_d3;
            oufl0_d5 <=  oufl0_d4;
            oufl0_d6 <=  oufl0_d5;
            oufl0_d7 <=  oufl0_d6;
            oufl0_d8 <=  oufl0_d7;
            oufl0_d9 <=  oufl0_d8;
            oufl0_d10 <=  oufl0_d9;
            oufl0_d11 <=  oufl0_d10;
            oufl0_d12 <=  oufl0_d11;
            oufl0_d13 <=  oufl0_d12;
            oufl0_d14 <=  oufl0_d13;
            oufl0_d15 <=  oufl0_d14;
            oufl0_d16 <=  oufl0_d15;
            oufl0_d17 <=  oufl0_d16;
            oufl0_d18 <=  oufl0_d17;
            oufl0_d19 <=  oufl0_d18;
            oufl0_d20 <=  oufl0_d19;
            oufl0_d21 <=  oufl0_d20;
            oufl0_d22 <=  oufl0_d21;
            oufl0_d23 <=  oufl0_d22;
            oufl0_d24 <=  oufl0_d23;
            oufl0_d25 <=  oufl0_d24;
            oufl0_d26 <=  oufl0_d25;
            oufl0_d27 <=  oufl0_d26;
            oufl0_d28 <=  oufl0_d27;
            oufl0_d29 <=  oufl0_d28;
            oufl0_d30 <=  oufl0_d29;
            oufl0_d31 <=  oufl0_d30;
            fixX0_d1 <=  fixX0;
            fixX_d1 <=  fixX;
            fixX_d2 <=  fixX_d1;
            fixX_d3 <=  fixX_d2;
            absK_d1 <=  absK;
            K_d1 <=  K;
            K_d2 <=  K_d1;
            K_d3 <=  K_d2;
            K_d4 <=  K_d3;
            K_d5 <=  K_d4;
            K_d6 <=  K_d5;
            K_d7 <=  K_d6;
            K_d8 <=  K_d7;
            K_d9 <=  K_d8;
            K_d10 <=  K_d9;
            K_d11 <=  K_d10;
            K_d12 <=  K_d11;
            K_d13 <=  K_d12;
            K_d14 <=  K_d13;
            K_d15 <=  K_d14;
            K_d16 <=  K_d15;
            K_d17 <=  K_d16;
            K_d18 <=  K_d17;
            K_d19 <=  K_d18;
            K_d20 <=  K_d19;
            K_d21 <=  K_d20;
            K_d22 <=  K_d21;
            K_d23 <=  K_d22;
            K_d24 <=  K_d23;
            K_d25 <=  K_d24;
            Z_d1 <=  Z;
            Z_d2 <=  Z_d1;
            Z_d3 <=  Z_d2;
            Z_d4 <=  Z_d3;
            Z_d5 <=  Z_d4;
            Z_d6 <=  Z_d5;
            Z_d7 <=  Z_d6;
            Z_d8 <=  Z_d7;
            Z_d9 <=  Z_d8;
            Z_d10 <=  Z_d9;
            Z_d11 <=  Z_d10;
            Zhigh_d1 <=  Zhigh;
            expA_d1 <=  expA;
            expA_d2 <=  expA_d1;
            expA_d3 <=  expA_d2;
            expA_d4 <=  expA_d3;
            expA_d5 <=  expA_d4;
            expA_d6 <=  expA_d5;
            expA_d7 <=  expA_d6;
            expA_d8 <=  expA_d7;
            expA_d9 <=  expA_d8;
            expA_d10 <=  expA_d9;
            expA_d11 <=  expA_d10;
            expA_d12 <=  expA_d11;
            expA_d13 <=  expA_d12;
            expA_d14 <=  expA_d13;
            expA_d15 <=  expA_d14;
            expA_d16 <=  expA_d15;
            expA_d17 <=  expA_d16;
            expA_d18 <=  expA_d17;
            expArounded_d1 <=  expArounded;
            expArounded_d2 <=  expArounded_d1;
            expArounded_d3 <=  expArounded_d2;
            expArounded_d4 <=  expArounded_d3;
            expArounded_d5 <=  expArounded_d4;
            expArounded_d6 <=  expArounded_d5;
            expArounded_d7 <=  expArounded_d6;
            expArounded_d8 <=  expArounded_d7;
            expArounded_d9 <=  expArounded_d8;
            expArounded_d10 <=  expArounded_d9;
           end if;
         end if;
      end process;
   Xexn <= X(wE+wFIn+2 downto wE+wFIn+1);
   XSign <= X(wE+wFIn);
   XexpField <= X(wE+wFIn-1 downto wFIn);
   Xfrac <= X(wFIn-1 downto 0);
   e0 <= conv_std_logic_vector(76, wE+2);  -- bias - (wF+g)
   shiftVal <= ("00" & XexpField) - e0; -- for a left shift
   -- underflow when input is shifted to zero (shiftval<0), in which case exp = 1
   resultWillBeOne <= shiftVal(wE+1);
   --  mantissa with implicit bit
   mXu <= "1" & Xfrac;
   -- Partial overflow/underflow detection
   ----------------Synchro barrier, entering cycle 1----------------
   oufl0 <= not shiftVal_d1(wE+1) when shiftVal_d1(wE downto 0) >= conv_std_logic_vector(58, wE+1) else '0';
   ---------------- cycle 0----------------
   shiftValIn <= shiftVal(5 downto 0);
   mantissa_shift: LeftShifter_48_by_max_58_uid41  -- pipelineDepth=2 maxInDelay=2.642e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                rst  => rst,
                 R => fixX0,
                 S => shiftValIn,
                 X => mXu);
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------

	-------ADA:MODIF'
		Tmp  <=  (58 downto 0 => not(resultWillBeOne_d3));
fixX <=  fixX0_d1(105 downto 47) and Tmp;
   --fixX <=  fixX0_d1(105 downto 47) and (58 downto 0 => not(resultWillBeOne_d3));
	-------ADA:MODIF'

   xMulIn <=  fixX(57 downto 48); -- truncation, error 2^-3
   mulInvLog2: FixRealKCM_M3_6_0_1_log_2_unsigned  -- pipelineDepth=1 maxInDelay=1.48992e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 R => absK,
                 X => xMulIn);
   ----------------Synchro barrier, entering cycle 4----------------
   ----------------Synchro barrier, entering cycle 5----------------
   minusAbsK <= (8 downto 0 => '0') - ('0' & absK_d1);
   K <= minusAbsK when  XSign_d5='1'   else ('0' & absK_d1);
   ---------------- cycle 4----------------
   mulLog2: FixRealKCM_0_7_M51_log_2_unsigned  -- pipelineDepth=2 maxInDelay=1.82472e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 R => absKLog2,
                 X => absK);
   ----------------Synchro barrier, entering cycle 6----------------
   subOp1 <= fixX_d3(50 downto 0) when XSign_d6='0' else not (fixX_d3(50 downto 0));
   subOp2 <= absKLog2(50 downto 0) when XSign_d6='1' else not (absKLog2(50 downto 0));
   theYAdder: IntAdder_51_f484_uid61  -- pipelineDepth=3 maxInDelay=2.03444e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 Cin => '1',
                 R => Y,
                 X => subOp1,
                 Y => subOp2);

   ----------------Synchro barrier, entering cycle 9----------------
   -- Now compute the exp of this fixed-point value
   Addr1 <= Y(50 downto 42);
   Z <= Y(41 downto 0);
   Zhigh <= Z(41 downto 9);
   table: firstExpTable_9_52  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 X => Addr1,
                 Y => expA);
   ----------------Synchro barrier, entering cycle 10----------------
-- signal delay at BRAM output = 1.75e-09
   poly: FunctionEvaluator_68  -- pipelineDepth=10 maxInDelay=2.19472e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 R_old => expZmZm1_0_old,
                 R => expZmZm1_0,
                 X => Zhigh_d1);
   ----------------Synchro barrier, entering cycle 20----------------
   expZmZm1 <= expZmZm1_0(33 downto 0); 
   -- Computing Z + (exp(Z)-1-Z)
   expZminus1X <= '0' & Z_d11;
   expZminus1Y <= (42 downto 34 => '0') & expZmZm1 ;
   Adder_expZminus1: IntAdder_43_f400_uid107  -- pipelineDepth=2 maxInDelay=1.96372e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 Cin =>  '0' ,
                 R => expZminus1,
                 X => expZminus1X,
                 Y => expZminus1Y);
   ----------------Synchro barrier, entering cycle 22----------------
   -- Truncating expA to the same accuracy as expZminus1
   ---------------- cycle 10----------------
   Adder_expArounded0: IntAdder_43_f400_uid113  -- pipelineDepth=2 maxInDelay=2.186e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 Cin =>  '1' ,
                 R => expArounded0,
                 X => expA(51 downto 9),
                 Y => "0000000000000000000000000000000000000000000");
   ----------------Synchro barrier, entering cycle 12----------------
   expArounded <= expArounded0(42 downto 1);
   ----------------Synchro barrier, entering cycle 22----------------
   TheLowerProduct: IntMultiplier_42_43_unsigned_uid119  -- pipelineDepth=6 maxInDelay=1.127e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 R => lowerProduct,
                 X => expArounded_d10,
                 Y => expZminus1);

   ----------------Synchro barrier, entering cycle 28----------------
   -- Final addition -- the product MSB bit weight is -k+2 = -7
   extendedLowerProduct <= ((51 downto 44 => '0') & lowerProduct(84 downto 41));
   TheFinalAdder: IntAdder_52_f400_uid133  -- pipelineDepth=2 maxInDelay=1.87172e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 Cin => '0',
                 R => expY,
                 X => expA_d18,
                 Y => extendedLowerProduct);

   ----------------Synchro barrier, entering cycle 30----------------
   needNoNorm <= expY(51);
   -- Rounding: all this should consume one row of LUTs
   preRoundBiasSig <= conv_std_logic_vector(127, wE+2)  & expY(50 downto 4) when needNoNorm = '1'
      else conv_std_logic_vector(126, wE+2)  & expY(49 downto 3) ;
   roundBit <= expY(3)  when needNoNorm = '1'    else expY(2) ;
   roundNormAddend <= K_d25(8) & K_d25 & (46 downto 1 => '0') & roundBit;
   roundedExpSigOperandAdder: IntAdder_57_f400_uid139  -- pipelineDepth=2 maxInDelay=2.36176e-09
      port map ( clk  => clk,
                 Enable => Enable,
-- OL                 rst  => rst,
                 Cin => '0',
                 R => roundedExpSigRes,
                 X => preRoundBiasSig,
                 Y => roundNormAddend);

   ----------------Synchro barrier, entering cycle 32----------------
   -- delay at adder output is 1.013e-09
   roundedExpSig <= roundedExpSigRes when Xexn_d32="01" else  "000" & (wE-2 downto 0 => '1') & (wF-1 downto 0 => '0');
   ofl1 <= not XSign_d32 and oufl0_d31 and (not Xexn_d32(1) and Xexn_d32(0)); -- input positive, normal,  very large
   ofl2 <= not XSign_d32 and (roundedExpSig(wE+wF) and not roundedExpSig(wE+wF+1)) and (not Xexn_d32(1) and Xexn_d32(0)); -- input positive, normal, overflowed
   ofl3 <= not XSign_d32 and Xexn_d32(1) and not Xexn_d32(0);  -- input was -infty
   ofl <= ofl1 or ofl2 or ofl3;
   ufl1 <= (roundedExpSig(wE+wF) and roundedExpSig(wE+wF+1))  and (not Xexn_d32(1) and Xexn_d32(0)); -- input normal
   ufl2 <= XSign_d32 and Xexn_d32(1) and not Xexn_d32(0);  -- input was -infty
   ufl3 <= XSign_d32 and oufl0_d31  and (not Xexn_d32(1) and Xexn_d32(0)); -- input negative, normal,  very large
   ufl <= ufl1 or ufl2 or ufl3;
   Rexn <= "11" when Xexn_d32 = "11"
      else "10" when ofl='1'
      else "00" when ufl='1'
      else "01";
   R <= Rexn & '0' & roundedExpSig(54 downto 0);
end architecture;
